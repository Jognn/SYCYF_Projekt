��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&��n?��1ů��> K�-� �&�T�Ek/ֆ�\�놭5�DꢘP���+L+X�4��J��#�0�8���������l��jT��+�(���������6�MC!D�;�m�퓊D@v_p��䙋ⲝ��C_�6�Ռ��#�� ���	RD�4D��畓7���vn�H���0���fX����4 �CS�C`{��;�L����li��� y+����FD�p"��]���y��R��K�({� .؜M�������	^5���ɋ��&���&�@*���
e�� �t+���
_6��O<��7f�M��u���m(MrN����z�jL���@T`��M3��c�uQ�Y���%�dD���,�~^���y@Ga��(����C����	��G�86�S$��ɳT�ز8���:r��/y�[ݦڍ#A�����i�&<nU��<[5)�Z�-Ĭv���0t���d���"_���:�'-��d��*��q����_d�y�N-��~";#��������Y��؆���	6ZJnԷW��έ$Y�K�?�4���L�w�Wmiɶ��Y�?jx#*�i���F�m�E����O6T>]i�_�9;�!(��kH7�OS��_��[-M�((��lO�s�$�g�x7`��ZV�E���F��,9�j	@���]}<�ahb5~ãdl&I^�	v����-�@�@���	��!��d��`j[Q��� r��;f�i�.�m+UH7��/OV��c��������l��i��M��*'��?���G� SK�M��H?�מqT'J,!A�h���'� D��G�T�>��tw�ܻ��l.pRu\7�V-�T�V���CS@�ewf���H�*�cwl�H��ϋ��#�`IY�k����_��U�A#���z\�yz�~�cٽ�bl����S�&+s#�V��%��ӧ'A�N��qT�7a�t��$d��]sH8�G�?����i��i6�ˋKl<�O/���	w�C��:�D��]�l9�ތ�G6���Ccyg9m��<%���o�m:|0�\)!�)�2�*�y�e�M��%����� w�Y�.���,���E�ٗ��N�*��O�zP�i8:³��v�\ݏ*�P�?���`�l��F-U=7�g���w��ȩ��$���"5��!������{Kh��������k�$V,[No�"a�K��H��c&W���Xu3ѳ����i�uI(of���p4<t�Xzf��4p-h��,����<��W%P�)�������c�%w]������"� �ۭ��9�[�Z_���K���N��� �{����Z�@���k}]�s�yR��݋}�k���/���7�&�<�V�0��dG�z}af��5#8��N1�M ��Tl}JĖ�B�	�}E�}�A�	K����D'�R�g��=	������+a������%s,^m�����Ԝ>�m�����?��/ ��#]>؊uN�\���0}�ڇ�T���cj~9�I/g�~0��1���'`p�4��w�:�)�W�M�^�p�r8�^�XO�>j�̫h��BZ�T:�x��z����p<xͿ`����u%�����HM��@\�(��'��b�#d�O��b�i� �SY�L�Z
�=,��H�G�tu�>��^<�Hv��o�z�@�(&\����F��Fq� s�SW�Gv��/������bE���9b�g3D
�'��}d��s�3�KZ�+J��#ӎ���<0}����@A�k%߽����ș39���G�Zx�D�\i�i��6g��y��C%��M���b�L�VU,��`q�Lv�x^m�b�g��$)$�.��诒c!���x�!�n�s:�ս��"����R��d\F�w/>O4xY|q�Rure���&����>��A�%�+:b$��2ji���i#@����� FhBo]47�� �Ϟ�z��P���M���U�zai>�B�CQނ����&�qə�AD�i��N��'c�]��!���򀋂��A*j����Q�@�]���k��K�
K����K��Di���àM8-ю_	�Ç�~��
dt�����z\]�y��q��9��1����'�N����g2Ly8��x=W�EK8B{ʭE�s춦S�6�(�����;����{���ׁ�������0�޾�>�%�4�}䢸Bu�Z=�?���۸�hl��Ԧ+��Y҂+\�~̷�Eׂ�)�~�N�S�*F�98gzxĖ�M�s���2��F�f%����z�J�uWZb��vS���(f�>����-\1-7GLl�2�f#j�xv^P�S���BG�;R�P).䑄!��l�Q76�M1ٍ�,y��U����=7�|�^��?R�,b����Z��x���~ߎl�',`s��ç��eS9i:�u7u�.�2=�$���`­��J ��-crF�n��W �����*	D��a���:�Ef #��$�gwd��+���$�[���Zo��qO��[I��f��szh�p��۹� &w�����[j3����;IO���˄�P��o_����Dؘ=2�[y����2�mN���1�;�!������<�@���>0���;Jg�?����F�6�?͇N���s���Ó�R�0"�$��:�c4D�ע'dV���=��T��8{��b��t�=�ꝅe���D!O��F��4]��e�7�HMi5�a�A舯�����'���m.��u@���������N1H� ��?M�l�/G(
�:e䇁�cH��!F)��O����ǃ#�SU��t*�f^ᚎb��M�1\�{�T
:+�ĺ���J�F��rdԆR#�U�2�@1Y��V-SƖ��J��^yl�*	���q��ׅ!��_�@����E�5 ٍ�� `�q[����|J&{M��2R����&.86;ǏX���6��(&��7�F��T�'�l�zRpnaLJO��:6;����κ�S���W�����d�JP՝��H"���i��4�e'p왚Ke@�t*����塘cS�~���UI���nE$�v�0b�p�Jew���z�a�!�7�*����N���D��"�pL��Q�E���1��^а����ݡ=E�lSJ��
%�*٥�����U�u�)!�⾁�vS=+-Ы���#��c��xԣz�V�c�����]���^v����#�ӷĊf��
$�D4��fe��/�Ȧ 5��L6�[E4�ѧ��'�H�A�ڣ�e�&�K��oH��1����\���P=2x�U�)��� a�qF�D/��
M��p�#����x�QM�s�'f�:���#|{���@2���g�EF�Xxߌ�`�; ��ݝE�yY�Q����8�o}o�\���1���n�5��֜�̹ &��6;�O��x hg=���Cb����jَ��Cɪ�%�p�Ɖ�-�z��tN��0X � ��x�ob\�Ԙ2V\Al- ̑��?mD-y2�?`G��"����	ݑ0���ؘ�Ln��?�P�}���g[�L�0�d�v>�1J5b�d��1��lߊ���M~]k�Y�*�I<=�sWb����"�Ap�
� g�G��J�|��Tm	S݂Ҥ���F26�VJX��Iݺ)e�|�4�#~��<�����_Qt��e��^�������9��>Cr��t���u𦋽�%J�Ʋ���t����v��]:�154Wv��VS�I���6-ȃ6Hh֌�gl�A�o@�N�oȷS������$���5�N�V�-�x���&]��9��X����Nܪ�h6	xĩ�/�XmTf�E��5[I#}���Ƌ��;ܼh����?����yy��v���Ɂ>��.A���]�F����ض%�,����?r�x��6��ILXqi喍�n�W��a�)���r��]X���yr""�@��	ab}�������eX4��d�~f�6�7[��Sd�@��i.������+�I$=�1m��}��V��U��!m)t�n;S3��pܾ[)ыa���N���3 ���( �֌T@��!<�xt#�cv�%�lr��W+n��gmd�bB��U%g�;V\��?'6�e9:u�RMT�o�
��R����K+ȹmH����4�~�t�����Hѫ��k�(/	��/�e��J����|��u�N!R�C�J�",n0͜p�8� -�*e<O�X)C*>C%�!����Y�n7ع�,��*�:IC�.��0�o������M��\��#�\�qr��es���|f�o�,X�o����-�8gn�ً0��g�;5K�;ٹ�>�Fu�'◷���������� U��t��m�<�@J7�h[�E�E��Ǯ��F�Q����	<H������щ��<1_o����g!������Ԣ��p..	[���EU�Y�����,>J�]�O'�|�۞X���TSPsO�.$��m�����;���D%�1�� Ői��C���%6�x�oDSi�_y����xk�����_��31&*1x]$U����:�9��Q*�[����|0����9�G5�w���Ʋ[�lc���0���b��p(�Z� o�b��[��
9�� ��-��Dz����!�?R��n`}�'!T�>�[���8�����5EG7�?5s�O�Xx��c��؄p�]���xݠڢ"r��	k�0�b���s�TQ=�а�e�<tז?�)OEr�.i�X��)�/�,_�	����nCP��Q�6������ud �}��; �H{~�כ�`7�SK��l��"�xb�fHHR�@;SjS����W��.P�y2WS��o��.�x��,���e'2V��ͱ��v��]耻�윝Te�=���gEu}�*]Vױ��4 ���_��nXY��8�3Y}�ٮ�ANj� =��3#��V�����S.l^����H�Jg#�b@��8<�\���[r��;2�`�(t.�R�q{�`�H58J��x8�Nm{:lli�;�9M�|m65|$�ۨ��G9Ѿ
��F	�w4ۿ ,').�[���K���pV7���
���I: �)�m�>��|��6�p�S���ШᲴ�j��M���_(��[��F��hj�o��j�;C������W<�0uؖ�靱U&Ag-D¬R�g�3��!�ib�#�ut�2&Ky���9.1�3SQ'f�3#���&H���3b���N��C���A:%{u)�5W�^��	�ܖ9/~�N㉂%irETf0�0����Ԇ�c�S�XsWl���I5 .q�f聽���xd�}��Aཛ�n;ǩ��L�̸$�h����AZ?��A�1=hk�N��Jn�4���/������6���P�"w�2�҇��&y��@2��e	V%6�^jh󻒺a�XX����Z% �F��Ν�>��X ����� Nԫ޸$�`�''��_��n�&Y;5R��z��A�����Q4e#�}U饳+�@FV�<�a�F tcQ�@\����%tv&�zα���W�l�ˌ��A^�O*��ц���r�2������P^���[iz�Y��}E��T ;����:VFH�_n��_Ÿ�� u�y���+�ݼk�����G��%'	��u���3�H�� S��9{ì�2	:�����fX�����|�Lq�.��� ����>¹p��0T""���X�Q�-n p)B�fS^f�G��ȷ5ee?Jap��}��;�o��D$S˅2���!�)���� ��,Ɲru��v`M��:4t����\I|�[�q���^�gݚ���n�9l�Sc����Ɩ��57�m�3�G�g�]p�[G��F;��z�O���x�qoG+����(�P�>���E�Y��S���魦�H>�>�1�y�!ʦ㌙��PO�d�8K�gۄQ�� �EWw��Ɠ�F��5#Z�W֯����'5߯Z��Π*h}�@pJ��$b��XLVn���1�~��!m
�>�^6Ӳ�NF���,�q�h�
IЗ���J�рV�Z^V/li)-���;(v׉��r��8��T#�!��g>ڠ&�}�D�����}c���f@]w��Q����r��O��̈́��l�'Rz��C�h"�տ�����zC*�y�
�fg�;w�՝��M�ʭ��(>WK�APs�u�D��E�D�Z�y�>�b=�]�gr��\��+���i/}Y�(;�)��_��R/'���H�=^�C= �σ�IY�q5j�u,�'|T"������~���7z ��*P�a.����`/��D��P7c��FO�+�#�jm�X���|u�e�x�ߒ�_O�VxZ9�a@�􃌼|���#�#w9�t�3�������֡����,PN�PȖ�ٓ��Ry?�h���D��OJWT;��Dt,
yL,�`e�$p��c}w���r�T�S.�Sw88j >��
+9���k��P��v���z��P����3]m1@S*L��`��9�,�չp����=&Z��r��.P��xIC���D��_��{�8@��8����&��}u���`}�8�{�HrG���%�ծ��uC=k�(����l��(��6��s�T�վ��	k�CԩQh7_PJ�d���k��Z�<��@d�t��w��`^}P,�L)����J�f�y:4z�齤��1���.���O��	�ΗTg�_i�x���=�[�ݛ�霊ܩƗ�KNVǍ$۷I��[o�Ƣ/|,^����w�����vjpm( ��Gx�Hښ���,���J��x�Gtı�ߣ*�k1~p��V�����;��t�g֯;�������a���H�����K9I�$�1݇����1�D�f�N���hꁽ]</Y �����r�fd`c�,���̧QRNbd�n/�0��� kA�%]_������{���L��ʏ�h����7��9��D��A�12��I�+���;�����N��o*�]2&;յL,�N������v��$9�My���U24���eJ��@1������3RDb��8�s��(w�7�2ֹ������~x�r���xd<����Ǜ�F��r ���F�p�`��{Hu��t������71G|z��'�	�����K���_.kh�R�����KH�G�����J ��-)��ճ�)�
ʥ���\�	�Yʽ__A�	�n-�
G�7��}��*� �^�ŏ���2Hl��{A�CV@!4�Y�=���F�d�N��߼(�����y�{�'15��i�CR��4X�h-�~�Bi��i��IW�\�W����4?��R\�e��/�������T�Ac@?W��;i��=��'�.�L����S=G���S�D�N����d���X��6��6qMv[*�E.�v졀zk.�p��y�F���2��+���6�Ϫ�0�<CZ������5@]��OG
g���`�p��e��X�ҚYJi�+�T!�C��g\p���o�)"Z����%�ڼގ~�(��'l2�0���
>��#6{[��.*����u�h��)�r�uT|�E���f�p�T���^���1�cH�ts�d�c���)������S����#e�O�wߓ��y0{YQ���mD��]�6 Di5�z6�:y�XV������v�]_�����̺N9�'ے��l�f}�js��\�h���,M��a'�c��u�[fB�jkڰi�oY�-%��.8A3�"���m����HH��a=��?ge�OPv�Ho��D���'���T�o��T�x�AN�|�v��࿔G�/�*�p���!��5�� ��-AH��Yso�I��	��)8`pR����q�*��� �l�{i`��D��5�O#H�����-�����f��*ѷ���㮧c`�g