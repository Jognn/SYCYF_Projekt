��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&��n?��1ů��> K�-� �&�T�Ek/ֆ�\�놭5�DꢘP���+L+X�4��J��#�0�8���������l��jT��+�(���������6�MC!D�;�m�퓊D@v_p��䙋ⲝ��C_�6�Ռ��#�� ���	RD�4D��畓7���vn�H���0���fX����4 �CS�C`{��;�L����li��� y+����FD�p"��]���y��R��K�({� .؜M�������	^5���ɋ��&���&�@*���
e�� �t+���
_6��O<��7f�M��u���m(MrN����z�jL���@T`��M3��c�uQ�Y���%�dD���,�~^���y@Ga��(����C����	��G�86�S$��ɳT�ز8���:r��/y�[ݦڍ#A�����i�&<nU��<[5)�Z�-Ĭv���0t���d���"_���:�'-��d��*��q����_d�y�N-��~";#��������Y��؆���	6ZJnԷW��έ$Y�K�?�4���L�w�Wmiɶ��Y�?jx#*�i���F�m�E����O6T>]i�_�9;�!(��kH7�OS��_��[-M�((��lO�s�$�g�x7`��ZV�E���F��,9�j	@���]}<�ahb5~ãdl&I^�	v����-�@�@���	��!��d��`j[Q��� r��;f�i�.�m+UH7��/OV��c��������l��i��M��*'��?���G� SK���mkݛq�K� xwC��f*CU+`�>�zkS}>�����{���K3�&�4�N�����Nؤ	$̂lUPo��t�-ME�U��j�Ì/����$��_s*���j�^��<��
�ZJ�S����C�N��,�J�e��$,%�Z���i�>�B�i�1~X*�P�}�.W95�f1�t�~�)��³O`��P�d�n�������P+��5�@��ʝ���80�ꬵ5Ϊ�յ9���މ�qR��q� ��� 3(�܏P�U��ŀ�i&k�⑭{�*��+E�$+��Ei~ܮs�4���Sb�� *�[-��hj��y3ƕw7� �<�XV�=�%b��d�Iy97�������c�>�^P�m<��H��8��ȇ(lO�Si:�m��}*�����g/��[�m����G��@9�M�)dl#���_Ρa�akD"|�Z�[��OT?�2�yʁ.�M���=��|�O���jJ �	ڼ7�(�PV��2��s����gWjw�P �|�Dc���R
߲f��%]�2Oor�Zc�:{͑�iV�|��H�쪤�L=�}`Х���&�r;۪��7�0���CB��i�>�)_��T���to����'v�nB�	I��q��$. ���,�<*|p'O%�1�����֦�?���)��6��L�b�� 5�m��/�D�Taло�X�<G��%S�Nd�MӁ�L%X܅Ŏ�F�
ܒ�#���RɻvJ�Ǣ#��y��e��uWs��V���%���CЄ����1�qp7J�_n!#|�b(����˺2��@X�����g���Aެ���@�~IG��$F�Ǔ��x�4�G�tR���g���ӊ3����� $�k
�e���cCj�0=�T��'D��d���UF*�+��~�����87-2��0( ]no�~�b��6�'S�m��J��{��y�kY�<Cm6�L��Z2c
�[�SZQ�*u��q���ӚsYt�ǧ����.�,����eJ��3� :���9Q@��5U:��M�Ŀ;d���i�I�]�<qnڭ9���`�p%��|��s�}�{s��7��^��f�Oƍ�]��M����bl~�l���UV��:�!���m��j��;o%���9h+�b�P�M�g�"6�|��l����f����Z��_��3��1}��%��|�@(�O��X�R��{�F;�� ��Hl��#�?������}6ɱ2#��!�\�0�K.���F�yx�&�8K#z���#zǇK�'�PO�/�~결�nͩb��`�n��Y�d�	�C����nO�UgL25l;��>u�y]���.��~�<k�]9�9󀳁�Z'�~]��虘A���3B�*���3�;�g���W�R��O��B]$b1�x>�g6�ԥ�����	6(/�s}ƙ�H�7䣹�)=+�]�E�f���i���G�oCv�ȿ��7��56l��?5�9�	�I�ټu%pqjOI�=?��c�U0�?����>���̛�-�s���Q�qX�������=P�m�C��
�t�2|�U�Q��[f4��v�#
lCc6�b�;��FiPD@�뻮,�RH���[(M���G��G��)K�mwۜ�}���XosXmcY��3�q�"_�Zjlt��EӋ38�h0����km��D(�>���]��nd�c�k얀�1:��I7B��9���I�-GW*a�\���<*�K���!���b�R@ JtE��i�c��v��+C�3HZ�@\�v�7Wd������}_���z`�T�bg9o�W@���v3QI}v���@�� qDF�G���!���vq�*�:01���$+�O*Ҫ����t.�2�٧��zy�:���x=��]���=��O��V�C�[Hm����'���Z'��%q�cn�GR_����'�	q�&�_"?�������y�`qgF��`��8�����ė��ǑX��������II���+�v�?�G�=��ݴ�9����=�B؄7�5]@���o��rh���S6"�'���(����U��%��;'⪻f4�ŏCh+8��e�^����F���N@�C�
$��R��՘+  K&>P���#hlib-�E�֙G�D��q���7�%���]�B^5a���������'�0hNMH�W+y��`EEvl��^=�W|(O	�`�02���ӗ��B�HBd��L�n��c�S��Vӫ����
�C:8�*�q"+Wom���L'��`��"!�� M�C�D�����{P!Ʌ�Y��� k�*�IqX�� 4:�,+��r+�9K8�q�W��RR�E:Ǔw���`���6�<&�c:J_(�;�vJ������%e�sh�<d���:�X�7��7�#AO?���2"�v�AV�W��������hl�P���Ν�O<oV�X�S��W��Cқ����Uf�8����dB�kp�1�#������X]�T�F'%�T���%��ޒ��?;�	4��J�8ɣFh����_�cn���nH,���Z��U,;��'���p����!n$��!�P  l޵�Cbn����-�]�CWABݫ�����c{oN�/��V���$
Y#��h<QZ)�b���;�u?��!TW{|csm)�|V� ��(2*���ڡZ��'q#H�'��"zM��հ׷V��6�g�м�3��7W�<�qgCz�ÿ��)�c.�9��k俄��𕸢��z�0���n�C*<J�>�&Vt�����A����ײ:80lB�����ON��;��8�J}��=�&�;�l�浟{
��UljM�7/cc�TfL">�V����ٿi�j�m� U!��ˏן�.j�Y��c6�4^���ÔǦO�DB���R���9�f��%N:��2�S��o�
9&V`re�b6k=6<�q����Arr�B��1"8��gh�(1��ٹ��6� ��S����L��\�7�k�t���� �Z���C7t ���� ���_ug���T��5Eݏ5�vZ�έй�!a&O\,���x�\,��⻿�'�dW�YHM:Z"���O�=�}{ ADn5^��fゝ�&~���7s{SE|e��*�:����Pz�&S*�O��E?���F�0���� �.`� Q30#���'<Q�Ƽ����W���Ǝt��NO����K`��8FaJ�G.��FW�_*�p�܃�X]�/���u))H�-˝k�+-ּ^�����u#/�߃�2HF��S02�ز�1����~0I��0�q%�� ��ߗa/�UyW��B̸Z�J ��j!����4i	��j�����%��kraM��3�(�����O���3�@��,�R�35��$%�w����)�d�^�mIW)3�@�.g,�f(u�sJG�I��I�Kz�Bs��-�Gp���$۔��&����&in��>��em�]��Gg�U��/TK��w�ӼJ�3d$�1{Ir�����f��Q|Le�Ba�m��p	
�4�T��`��ߐ�_��F�[�h���Ku��vBo������6�}�6~��Fw� p�!�sy�����W�x��|䗃@\���=@�.X:FD{Q�G�����P�ڟ���["���`rǟ�B��s!���_�E���Ca�bb|�;��M��,s�n�k����-|�=�~N�ޅ^��ہvo��+���hAR?|�*l�v��)3l�#�WOa��9_�ȴ�HT��� ��L�����̌h��M��d����)ni«�	.�\Ńr|��2���>n	��X*&[�W�-�A���|�3)��;oUņ��m}e#�m�vq��~L�]3���O����.B��*e�!Z����D�O�Ǐ��i�'�������¼dqN�O_j|4�`2���4�Q'	���qD%�{�c�.�x�γ:��hp���N�['�� ��� {���F��<�vj)PP59ù�E����$�w��/�l^�,��!4_��M���;���S��_�J���p>KT�[$��YO�_�����縀c����Sou�&^��pX.�x�L^��K����^d��'�p�
�+��P���q6�v��.V{(q���H�H	���Sǫ8����}���X�b\��A~�˟d��Di��{�<�c9|T�yS���Y��U��i	�H�݈�W)�nz�=��_��IaI�D��u��]��k�k[ԩ҆0C�N�q�y�S7Q| ��dgӓ����]ߺ^�q��� \�JPXɃ�+���o-p�`jM�:(��?�܅n���o�:"�/$�R�F��]1�('D$��b
�U��Gqc�v�^I��:�_��r ������{�A���?w����@�)�;����UF�妬7�w�Q/~^m���$�ڜ���������1ʑR���KKF��@(h�ƹ79�D�+��n���;�-�<��+=!豃1w���*|4��#?���J �>|�`Ӕf��P�r��8XV�KdH�H��!8��*"��`J�O��Ě��DD`�W�%=����|��{%��^\<́��2u�B^g���wQO��{uh�b8m��MA����Oa�ظ?.�PWi(J2x�u*��n����{b(�Y� )m\�t߼v���Yө�*��%wІ�s�+�2b��|
 h���Q�q����9Et���<>Z�3��0q=�1Q	O��ڛ$Gf�����͟d�Jѻ�B��-����~|��2��p�0p�a��I���,ԁA�PL���ə	�K����k��خ�����]H6L�]��P�o��S>F��d�i�q�&�WM.��G��u��V�B�t�V7d�X���
��i�6&C�'~���b��Q-d�.���4��qGؚP�<!|�Q?���D��.�����1n�3��#���7����⤽�,q>���b��,) Th�q�����zP#;7��[�;ϭ]�f�%b���BZ�}�x�/sY�'��9�n��Q:uK�y���ŧ+�wFİ���b" �y�=M��I�F��T�܏��y9ڥ�D��� |,�l����~x
cB7a���_��C�P��('�,��\!�z��{7�|\c�$<�
(B}~JH����܎V����vr�d�c������a
�k��i9Ѵ��2��>E�A��R�o��Ȩ�
"	���#�Ύ���!�VAq{f�I2إ��<@�V)�B	�����t�R><�a7ywUDYO�'eV90��@�Y�P� ��Oǅ�R
;*C�HAn���@��f�VV�@��(�&���,�4�=���Q`�:\�����=���j��^Æ�V(�>��}��]��c8E�Hb�$
�lB� ���)�����(�%�y0�����f�
��"��XC^��_�Ov����3���E����	�Sλzw�U�I?��t1��U@�:vA��3b��mR<>�yB"X~"A����qm˴?�)�$M�U�gĵ�&�R��.�M��X$��G�|5���Y������3�=j��+�b:Ab�R�	av�(J���]�����%�� Y�Pd�=,�@H��'R��������aAL��7��0�m<~�]{�P"ɞ��0@�Z�>����mi5��̙��X�A�G���?��uŁs(Gm�ؔ�*�f��E�*��jǬ���0B%�ag,f�"��	-��ğ��⸞u��o��]7�M!15><�����:s�ˎ�:+�8CPZ$Ƅ��}�s4i��@��f����E��t�{6���7�%HV�iޗ��?��W�2O9�s�bD�^Ŷ夵|�nhN�V���tzH��E#��&m�R��2_Gs��U�9�N���jb-?X�K�����kK�|/��lR�9DI�]�ƎH��H�Z�t��_qNZ�V�?��I�I�]�i�%�~_��.&��lT:���F}�I�K�_��F�-�b��$��iX�x�����
�|����	��:��~�O� ���+�N���kA��z�o ��(�k�<|['��/nR.��c����]����G�$C��W̚EU��Z�	�nWtӜ�ϕ�|���H�5����:u��O	��<>R�<a��/���\��Bش�޺	���!�2�35�,X��lJ�+��U�{ �_J�b�U�����b!�u�%�Bk��*�?�$� .�Ӯ�7��}�j�^��&Rl�>A$�V6o����<�e�}�l�0P���.�-������S*��t��cۂ�v˅�}���I���6X�̂�l��=5(�Z��C+Y@������u�l������vd6��	��(��}e̶�r-���L�1�]�N�ߴ!�� A5#�X�����S�i��ʙ;N�R�a��z�X��B�y\�H���wǬ��O
�!��9-�=[5���>��\m�tk��_ֿ�#��=;I��_������x����%׵V��n6]��ٜ�m';��}ͯ?����9'��X��� p��-�]�6��.�a*v�����Y,��=�p#�l�*���a��t���46�?��IgpJb�u�E^�EdAa1�N�0��YG#7���໌8�.�T�E�m�>]̛�/�A�0C}�)��9�!��n���ϰ��G�%Γ�x�?~$:5�O�4~�s\ 6�*:�G�C ���i8&D���=pq����HS��1q��'�i]�3,	?CF̲�=�+٩�j)坋�0Q�8s�K���Նɦjza{�D# '��4�lGoGYPk�Č�l{�Pl<g~aJ�D/O
�o�<YP&8�^�䬂�d��U���