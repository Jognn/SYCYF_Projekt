��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&��n?��1ů��> K�-� �&�T�Ek/ֆ�\�놭5�DꢘP���+L+X�4��J��#�0�8���������l��jT��+�(���������6�MC!D�;�m�퓊D@v_p��䙋ⲝ��C_�6�Ռ��#�� ���	RD�4D��畓7���vn�H���0���fX����4 �CS�C`{��;�L����li��� y+����FD�p"��]���y��R��K�({� .؜M�������	^5���ɋ��&���&�@*���
e�� �t+���
_6��O<��7f�M��u���m(MrN����z�jL���@T`��M3��c�uQ�Y���%�dD���,�~^���y@Ga��(����C����	��G�86�S$��ɳT�ز8���:r��/y�[ݦڍ#A�����i�&<nU��<[5)�Z�-Ĭv���0t���d���"_���:�'-��d��*��q����_d�y�N-��~";#��������Y��؆���	6ZJnԷW��έ$Y�K�?�4���L�w�Wmiɶ��Y�?jx#*�i���F�m�E����O6T>]i�_�9;�!(��kH7�OS��_��[-M�((��lO�s�$�g�x7`��ZV�E���F��,9�j	@���]}<�ahb5~ãdl&I^�	v����-�@�@���	��!��d��`j[Q��� r��;f�i�.�m+UH7��/OV��c��������l��i��M��*'��?���G� SK�M��H?�ç��q;��)��Rȩ�"@���r��Ml>8!�S��L��EgeH]�8��>]GR=&���C��i�Za�z�,�F��h�q��^���wT�a���%�9�n��?~SИſ~�mu�OlIv�4'sT���/a��^��9��*��G�Fh�DM�_��CN�<�_Pg��O5��}s�%��m�o߫R���X�Q��	:����tգ@�����K�<m�|E�F�_�ʊ?M6�)�C�,��B@-�/�B�����89n��Lq�N>�~]��5�|��p�)Lٱ��iM9���A�<�*j���92�E�F����Jj�ӟ���Di*+HB�S1��V����Ε1Qr<�dIX���	"�=*>p��[W� ��yRAˠd�Q�&	�16Q��m:�B���W��,��}w)tԟ�B����S�h�~��]H�=ս>3�b�>��i|kD����\��iC����<�Ӕ����_��Kj8>���^W�!gȾ[>U�tCK��3&��h}�|fA��
���t��o�>rmt�R���m��S���_^��� `0�RhP\���T ����1D�g��C�~� ]��4�c�g�l��:����לn�e+�����0Mq�ժ��0"_(@2:h��<���q�Sg=�pr�_VɨEf�����|_f���J��au��#yJ�F#n)(v���X�C�u���.1;IS닔ˈ�|�N'�{�N����	�YZK��>ʉk�v�����i<�r߼�^@�<��i1���\|P�gx�ǯ'V��>�����o�K-"3��A��0wa���JBg��h�1����I����dծ��{d�{�W��]I����*頃q����B<*�_��Z�%}7��\�Ͽ����M���D��_ugcS1�d�)Kk�t��H�y��c��^*�����<W(���1���:�$Q��
d�G�h�zֈQI�eZiz�H2B���
�;5���%-�H����$(�u-�cd�k���']� À˛������p|N����T�E���&;��t'T��V!ow�[��+�$M�����_\�/,�� �d�Н��2V��7��ݯfu��.�����Ք�:���|��M\F��)?������W�t �ˇ�,G��w9���7/���C]i� '�N��i>�t��Sֈ �/����u�3���3x(�(g=5ju�y)(��@���Y��s��5@he�<V�t
pi�n0�fOr2�r���<bŒ^��{�5g_��'��N���u ��=s40�3�=��;�W�'��]s���'F	Z�,v�m"����u���P�ԅ���������X�.40�0h��8�(@
=r5���(d��@�a6C��[u�;�A�eQA��g �Ω4�l�*�6\����tJ1�gk��4C��[���)W�}���7�}���$����D���$>�����vSL����TЎ��^�=BrT�y�Dm�O���O>���#����D0a�v,Yel���� !����7CF��?b����z�tJ��Ʀ;�R��"��6XeEº%@N��OI�����K�{�?��\�f�Q�7@��5%G�^�4�va�5�N��\qwy��F(�[uj�Z��&���Y�~4)�"o$uh�G�� ����{���M2�d���-����&Q�:g�GHa���T����{�DsE�sc~p�,�0���Ҿ&�t��zY��^�����̩�lOƒ�(�Qj�"��u���|�0i�_vX��7ə�b����R�~�(k�4қ�4W�D�2�+@g¬o��E.�$G��(�W�E���0��G��n��rr��^*��r��	���n��H���V/����{IY�y���-Mv�O3g��E��7b�u3���x�(�h�|�h���HL^b����E���!QAqzy��AI�w�fG h?=1��Æ��8		��\`Đ��*#�u���WEMz��)�h�xGr�Ĉ�2n�z�qڃ�a�}�+5Oak�þ�����FO���$��>���G=�'x�BW1�Gv;i�����6�}�2r�T6�;k��3���z�SK#��fQ�w�ZqVj�u<%&i��|�Tׯ��u^.	�v�bD�Z�e6����T|`�14��nw�C���J���v��ԍ:���y��Í�ŨŹi�Cd.`�Zƨm|�i�J��0l�	(��nP�ۢ
g�����[]ا>!y�n~��T���6��`�~N�|%�[!�]����ӟ�Nw�x[�MFd�v�҂B���ӯ0x�^���n8���+���@��G1���m��������N��s�\4�/e�N!0l�<�Fd�b���\$�0� �M��G](����M���dE�%U�"��YxӐ��Ǭ�^v�(�Yo?�)��Q��+%0