��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&��n?��1ů��> K�-� �&�T�Ek/ֆ�\�놭5�DꢘP���+L+X�4��J��#�0�8���������l��jT��+�(���������6�MC!D�;�m�퓊D@v_p��䙋ⲝ��C_�6�Ռ��#�� ���	RD�4D��畓7���vn�H���0���fX����4 �CS�C`{��;�L����li��� y+����FD�p"��]���y��R��K�({� .؜M�������	^5���ɋ��&���&�@*���
e�� �t+���
_6��O<��7f�M��u���m(MrN����z�jL���@T`��M3��c�uQ�Y���%�dD���,�~^���y@Ga��(����C����	��G�86�S$��ɳT�ز8���:r��/y�[ݦڍ#A�����i�&<nU��<[5)�Z�-Ĭv���0t���d���"_���:�'-��d��*��q����_d�y�N-��~";#��������Y��؆���	6ZJnԷW��έ$Y�K�?�4���L�w�Wmiɶ��Y�?jx#*�i���F�m�E����O6T>]i�_�9;�!(��kH7�OS��_��[-M�((��lO�s�$�g�x7`��ZV�E���F��,9�j	@���]}<�ahb5~ãdl&I^�	v����-�@�@���	��!��d��`j[Q��� r��;f�i�.�m+UH7��/OV��c��������l��i��M��*'��?���G� SK�M��H?�ç��q;��)��Rȩ�"@���r��Ml>8!�S��L��EgeH]�8��>]GR=&���C��i�Za�z�,�F��h�q��^���wT�a���%�9�n��?~SИſ~�mu�OlIv�4'sT���/a��^��9��*��G�Fh�DM�_��CN�<�_Pg��O5��}s�%��m�o߫R���X�Q?��dK�Z|:�=��y�P�)�� �\�-��d��jj����j�f���L��[N�����lhtI�Ĺ���ʗI��	��&P+��795Я��K��
�H�}g�G��ݧ�nD��t����r{��Q=�ξ�_����qw�APy�e�u�D�>���$'��)k���7����T4:1�ybi!�N������kX>]+�VFR�f{�m�*^���� #��n��ǳ+{e����r2gȏ�[V&�!�-�`yK��#�tO���=������ޏ�0u����m��!�F�GXI��H�6��������ɐ�=aPfߝ���V�xhw�\m&�����	�0��H�{�ڃZ0�N��w���/@+qL��=�|��W��|�R��kv�d��Gm)gn�茩a��ڨK�;uY.G�1Л���u�v����!ʹ���s�Wc�D.�|dE��J -WKH�g���f+����Ny{c岭�\��|�+�2��M��#Jģ�(J��2Z9�**j�-5j�@�鋉��nRC��͉��8�r]��fl��7q7;8}���k�ɣN����G���l��q�l�[�����d���V�{r�p1�,�ֿ�c3��`]e^������z�ܬ{+S�i�Q7�߶v|nQ(��ģ�_�l~�d%�$$���FB�Y��6_˱��#��6��J:��hl��p����Ø�p��->��d���U���;�,�	Ø%�L��|k�}u&�(ຜN�=�?�p�3X�~�����]��i��&G�5��[o���N/��n�놻�#�a6�E"�"wۤ�ǜ"O=Aq��-XV���\��I�0<��9��b�� aO���JC��d ��/�֌TYC�nGr6�OᯙI�o�Ϝt\�6�8AO�~��%�a<�.�m�E�:��bO��xC��7�t�"M������O��t,�iR��w<0e��`��͉��A�J��)j����^/�W��N2&��#�����i�l*�/�yhw�g�ϭ��9oy���ؾm�_�p4�cTX���x0_��`(xo��_�G��PĒ�y��)��ο�}Y>$���u��P>�<S�A΂8��(5i�6Cϐ���7�E.f1(N�i�� �¸�����U�b^�2�a�t|M��d�#�-�ů5 ��^���ۻ�y&2�Gb�F�f�w �y����~��n%"�L�ܾ=n�WP��O��d�
���� �D���d�3�F�  ^wUE��nz5B8`sp0$Kcn*��w�jG�FZ�e~�*���^�<�)�y�d8���A
*�k;l�E|��X����WE��@M:A���]���{l�EK�A��{0��ج��܆���.�UJcG�^
^�FK���{��-��!�"
���#�WR�_��os�Xl��a����D@H�ˉ)���I I�Є��B�8��nXRxns����S���«��;�����v��ҽ�������ʮx,��0|�m�;y!'��t��а���>BA��=��Pr
 }M�� ������O��( c�Ȳl�Dǅ�"��"]+K%�
�"����&^G��}�,�ȣ�k�'Q �H1m_�-��/N�]Ƭ�eI����e��k���3����Y�E}���M�
�6�`oFo+WakL��KX�����$�:u���X&c+f�\���"�2��P��F�x���'ӏ��BE������]Ȣ*9/�@ �1�w��$��t��#�M|�=�3�47��� �߁v�XwT��?��ueJ�'���1�FJ�>���F:jl��z},9Y4����� rJ����l
ղ"U))�$Hs���1��??!1W��RN�\���?�_�f �0��6��رd��f�U�h֝��~$�e����v�*��yz��PF{���&C¤(g%����W��Yj�+��y����|�,r�P�_�[J�ɪ�'(m�K��mԍ�#���4��)��~g$;�"�/?��3��*9</�%�9`����U0NޫR��_�_��	_'�s��������Vb�"⅘��EA�Q���V%�㥹 *@���E34,�z�06sR��A����A����mBe�;���J= �8UM��V��3�^Sk����/�j���Ų��3Ō^��Ӧ����ց��u�[��?>F��*|a<�9�|����b�:�K&��A�6{q�k.���\ݻT�������P���(�܅kOL��"�p�3��y@�-�v����xš9���ҍX�x��hhF��4=,��W��*
D�ٮwc�	bT1I��=1��V�n�˓�����u���M�Y=:'�PIG��g�3Fi����R��H�8�`��|��eE<֨�Q$Ҽ��+�Ĝ$��i�"���"��Y �����x�&s0���\���,_�C�f��L1�����r��3��.n�hNԆ�n�ep���[�H� Hu�ҢD
`������~�t�H���N�#�h�(P��9X�R���b����0 .f�;ґ�ƱG0$�H���'����`L��\W�S�OȃA)��H�Yv�ܡ� :�����B���Wv�C]ȃX�&��,�4]u��}Y�E�T�����M�X��w�J������t_t(�
)!��?�}LXףŠ!�4�5*wt��r�M*�+���*��1\Eb��!����^}6���t�����jsBV������z��\RT�Ur0�o����߈���d�>!�{7�Sϥ�j��ܷ��A݌+{�8������jO�NALǴC.!�N�a^�
`�I~(�g�
!�(K������9��jP�!�����~�T���S +�)�8�K��,���&�� �Z�*>�<�������]��/ڤ[�K�HGAw�s��E����I��g�TEa��7�$WFYt��&�A�ύL8��cS�U$Z�0�9��(=�.��\F-�N�C�PD@�l#ƃ���������;�uJ�۱�؟��bG�Ʉ8���Z��Y��;���)#���-�Sz?K%2�yˀ��/.����\$ʒ������<nh�V�m#��o Y�]R��ȰP5��٭�xR*)�����g�y���z�Hҟ�Z�>v繕Bn5����C�o5AT�Q��צV6�V�K3�W
��&K�����$nɎ� �;`@8��W��:�=t?�r��s,��p�"mǥ�;l��/+�F`o��%�4������V�b�&��7B������f��!Ӟ�?D<V'���"�(1����^�p�?���UrT}�E�uVAї����u��FH9��B3��QR�W�ʦq���<#x�N���+��J����L ��Gb�I*�6J�z�]�y�E�Qp~�E`��ʊV��>a�{�`0>���v�n�>R˘9�gkY�M:Y:�e����ݦ�P�c�}�td���+��؄����i�>��f�~⫯l�X�T���i�ca�'9����(��d���]m�E֌��A7���U��+P�f�5�j���1y&��7���W׸����޽z���0�9E�io-1��фo��������������������+j'x+Q��fI/%bm��(T� f�Yi��2�)��Wj�{Y?�B!��HdiAk,���!�?�ӟpGo���F����1��*YW������:#�k6Uۤ��X�ߩ�i'tE�VTEi�F���W�Vf�P՞(d�fR���=&���ykr��s��3U�r�B7���IZ�"C�zu�'>D)��0�#�m�;c���ᢌ)����T�|�	Z������Zg��SĒ�5�r+�I���|�Q�dBh��@��ԙ�U|^���	�����U-%�e0cy�"4�o�-�j�� F����cWp�8�~��ZBl�T�@ ��������)��?9|�:~eUҝY��k���Z�}�m�.�ᯋz�i�;��*�0!�����^\�(���$����0fBVc�{cpA���h�i������V'�QpF��t�E�6�W��[%| �BN�B��T��u+�}���Q��:���84�F�.�)�F��g�7����G����%b�UN0���v���騯Py�^1]��=�6%{�FF��	^��e>��ٳ	��7#zǍ��鑜�N3Ӯ�bX:v���t�{����H�vkB�'���vcW�5����(^���B��k\f%�y֊�POX1���}N`����u��ئoP����Q�9�13�
Iwd����=��C\Lc�C���M��LdVc����U|@�tc
WR&:p|( �hu�(dI��ڂ�#惋�|�O��Z9��XG�;U��e�@��+��{��A4��.�Fg��0rY���U��"�pxye!�GP<1�t�9~	���=�>J�ʎqM��+����IbM�I���y	ق��9���]�y�������"�Lш�h�]J�!=���hmY 
ه����k#��lj�᪭�>G)�ʌ�ɧVY>�Q����A���K��W�Q��eFj�%0�,kK.M�&�xF&B%_�c4kyP���sc��a��m�m�)<��`���N�(�\��X�B����`q?c�%`�z��S�+�O}8�W�*|��O:"��hr��R�v����������_�W g�s��-�!�UZ�'.wMMۍh.ai��+x}ܫ�Dr�/����X��Joq u���w��g�e��Aj
v�yVba�:�x�b����B&S+��F�a�݊��M���g�C��J��|k:���)ɰ�ˍ���;�j�-�!�2ll>���V��;`��B�&��4�%�9sJ1�*!뀙IH���?E��h;K�B?�pV	L;9��p�)��XhW%?�F��+�������pI�\�k.H�ң���h�p����m�����~�������}UU)ۢ0*�D6��Gq���욆�^\L�S�4�M������g8@�s��裣F��o����y��'P[	2�N�0NsI��?�;�S41���4L�Y�W���,�4���x+��N�Z��9���:dG���?���W�8Vg�4��^$*��1��cn2�%{s_�B�+��e�%.Q����_
��O�����ΐ'ETp��Id�]ݰ%;��Iʋ��x<c��z�� �=�����h}k.�J=\�Ddk�$�դ(���B�b Q؛C��[z#����$��)��>�������Y�嗴�Zq�����%�Bs�f�]��.}������j���S�bf�5��ȗ�O~ל�憴f�x�{�/Ly`ƿ��Z|��Ų�	��Q()�mLKW  ���;����є����U1/$�-jgN�Ο��g@`AuF#�'�y8�&���Dh�Ѐ?ʪ��zl���vQ�'�/j2��)	��iu��(��G���_b�L 8��e�Q��\�Ur�VG@{fC9�5}�R��U2�!%��������&;ط�&V_^�>�S�<����UY��^�^m(�P�k�?`��X� �(�Y�?��~�t�=�>�S	t�3LY�Bx��t�(���j7%c}�[_d��֕�L!E�O�DG����z���_nP�\p�Y]�� �l�L~�f|-�����]~xRb�E<7g�ǺS��Z���SyL�Ik=��O�@�!MQ
�u�~��ܕa�����ׯ�p��:�(�5)ޭ�:a���*o+�@O��Od�)�B�2/��Tqˎ/D�@G�5��˃��ò��T!u�^���*<��Nw
k�?�L�ME	CaKTB�ٙJ
����-�����bLFn*�t�4��AKr�3͏��fv�n��(Z-���*� ����i�4;�M��pfYdn�<�~Sh{��g���7iԙZ2�fz�_\5��ZE�K��ޅxk�dNX2Ȓy/��!��+�3)���{�ejѓ~������%{8��V_�S,�$ɱ|F>�}ޮBq�չ�nK���i��XP�����_lu�x���p�	A��i޲�j贺�%o0��R�W�8���Eh�K��Nto�Ӌc�٫��RC�j���(u�O�c�MQ�	�[Hm�8���o���]�{��L���;�sq��_�U��Yt���A��<9Fa���h�z�Hs���5_^;���>u��&�_:��T���CpPp
�+�rx{�<���W �u�{��3���E����b�񵞲lz��j��+r�"*�]�p�ƟT�cY�!�qf��`Uk���F�:wo�~N}��c�]�f
h�gpe����lg����<��? � �!e��{�с�p�y6Na�Ȼ�����K����Ma�X������U��9�!��l_%pP����1�����VWy��f~��U�� I���L�*�p8`h{�:uͽ�Z(�-��/Z��-���l]z�ژ�I�WC[�fL��|�Y�����P�����\T�X
�����`����-cW����S �)�T:p�g9.��W�gmn�Q	�uuT�� 9LO�$Ìh�.|ii`��>��\��n�!v0�)�A����'��i�{"�������?Ԋ��/�)�[��z,��SZ^�3��y�P+#��7������IקP��F�I~��F�ȀK�]��f����A�ɝ]m��&��.~2X�̆=�=WJ�h�];4��)����� ��ɎU�$��)&��:�����NVI��#�M�w��e�	+�����&�|�L�*��/���`����T27s�pWݵa6��k�i;e���Ϸ[���}�0���c��E*����mPONM�˭mT�p��̅6�@�u8��X���r��tt���k�!*
���5(���s���V	Sm�v��j����}�N���ڥ�iy1w�_sD/>�mad���?%��p�f�U��?i�n��-xͽ���p�R��I����;��~���^����-���Vׁ �E H�_�_{7�s�V:�5vF�`y�C���W�駧�k�Y�F���齉1�Ľ��� *%|��E���ӜPUL�d����"�����Y���<5���,n��#�;kF�7s{.��=mc�^�X����f9`SY�K�'��G �^��e��j|�.ob��yd5=�D�sh�w��yE�R������N]eM��#{��	�mY�m�tS",-νΐc�)&��/
��^(�W�7����i�C�1{X�ƕ��͜�K�n�Vj_\�VD�� �/�p&ӿn-�qI9aB�����SR�U']ʦG�t��'o��,�:)�==�/�0s 5X"(�����+�69�H.��WX�'�mb��H	a_=�1�����������% ��;y��q(oL>�<CS�h�Ĩ�6S�"3�lt��w����g�YЏ�3��񳸪+���KJ�V����>��$��a���Qt��1^Q�=�� ���*tc{��H� D���
fa|	+�����4+���&���Mya�!��e9�x�
?g�T�kj�u�+�{	X-[ ������=w`_���&=��3Z�<Gl�����K�⪠~����&]m]r3H��3�hb+n�9ܚ��_�!ZΖ�_"�SWY�r�nht٬�G��W��?d3�����4uY�RUTz��{B�.�;yb�����Oܢ�I��MX3_X����� {|~��s��3��a���&�M���m�v6�@�h�kb/e��5<�|��F�<d]Pl�cf>�	q�k�*"�g�u�Ө�?'c�j��@��ԆK!9x�>/X��"��l��i�z�iqo�o������[{ف6'��"��[}����p!�l�R|�3��=��'���I9\��>�;<z�!2֦,��Y��^����6j4���]y��.Z�5`<��!24n��i݀5D��L$F��Qȹh2�� �^�߷� 3�Z�"ѡ�[�B�� ��ٶΰ�\�:���T��eNFI:l૽���=��:��}���'��<B�6��y]��>�&(A��h3,aqt�/�P�&L����6y3�4ʶ�p�����)��pzz�k��ߦX����(1#������,�[�!���)<y�}���l/YAX�:J0��L�T��;��Q��t|��{��w���?��a��������hqٙ�;8��2�S�<Fb0=�'3K2�y���J��)}�W|����?<��6��;��2sd�l?ˍ28x��|�;��躰x�-hKϐ�P�Y��(���L[c-�]��v��PKb��-o� k��|������`s,�E�Wkڿ�'�럊�wP4]PZ!�� �����ŀ9�O��騫�S}��DY�G�"#S����eRU�����Y֜O���"IP�E�f��2{��iY!�ud��+2,��� �u�J��]9�@����y}�Ր�aT���':V\�]�`<w����*b�ͻ�*C��7Z� ��G#����ܼR��݃]q��~�H`^9�Ԓ���n:�ۯ�����K%}Cܺ[w�5b�9�˘^# �5m��p����_��'�~4������=��-��#ڢ�־}uI� l��ӈLaneo�?��u��a˰�����M����i����k,�ŧ�xS~�"H&:7�]1���u���0_H���6?�Č%J�,��%�P:��'�8V��Iٙy�B�m�<-� 
�d8;q���'�|i^MF/2N~u"��#�mn�fR��\�Z1BV�C�Z����o+�ex�;���F[���:��'5��T�Z�*�q��;�i+�h���A?|x�"�l�h��z �y��-���J������+������H<�:�8�������� S��?B^*g���u�Y{��5�A1���b�8ȡ��K��͖`�T\��"ثyi�8S=i��&�}���+&�V�3���f3j��Y+�*���<�}���v}$�j�D	zP��4q���C��{�T�������yƼ߲l���u�T��)_7��W��SH�䈉��5�r�P���m�j �RKb����%>��6��>!��$��T%�ۇ(\���O+�b�A��딍ga���Q-h9��s�A>R���8v�vD^��v���Pt��w�f ͧH���zW���*`� �5�wW1fŏ�?�<ƥ0�
�q���I��E�\u�g�z�K��,��6R��6n�U�z~�?�7�W!�|�����TEc��C�5�/�l&��|n՚�;/�����c���N����A�$QA ��D�L�/���*ÊX������F�U�iil�v<�y=�3Y�@�m���8�'8�F�SN���+��j�s`��~j�+TB�X���ɰ�ыί�U�D�u�Q�҂G�c(%7�:�8����yd撘p5�z�& QIL�@�����Ӛ>�wĻj�r4�"�n��H��ɕ.Pg⊰cP��|��:6Kc`S^f�+�c�A�ZȘ �f��]�s.J���m�EȻ@�
�8y��* .�?rf���
��ʢf�k
oN�=��l�˻-:��dP`.0m
���{!�4�����AS4@�Լ\��'t��"ԍ��1��Ŧm�U o��&�W#��'5yp�3��4I�^��:~�ƒ���sq��ۮ�ä]�d�A��.���U���q{Uri
wA|�D���Z�=�"P��3�ϸ�a�F�OÌ���Z��>��4�MB������RD��{�}k�=�����vYdΚ��	���s��mll`5E^�ϪU������\
���Y+%��2.��2�H������������@N1
�X+�$̢�{�j6A^ߓ�T���"gE�)�L�z�}�k�kk��W��rc��4�4X��� A�y�un�4GΑAظvI���:-_������ÅVl��x]f(��:����p˨v�e$H���N@���`U��?�7�"c��p��N�5�������f�G��es�MBw=������+ppjv�Ěyp�8h�s$�Ȭ��\LUjȚ�U�{�-'���]J�aZ� ��i0{�2�7�T%iD�I���%thϋ*SH�6���1�g��B��5Tz�}�3���Z��������o�)Ax$e�B�׳�j_�&tc�N�67;X	F��2�T)wv�@Y���5${lC#d��� o_s1��7���]��k�F�-"'�Ӓ=�bm�kg6G#����fS���=�/��O	���h�l	*Oԫ3����S:������
HH�%�
��wg����%��c^�@���WT�7�����HWGM��y8���T�3����ά��N#� i��� �`#�7.�%(�jD�[�}�.\�m����M�P��/������}��O�(Ը׀�(�\�O;rͯ�E�h>�~06��￠G���D&�1{:�*/���H2ԛ��)�d��8l��:���UEm�(�~:�PU]n{�@�����T�$��E��O��`�#��iE��|&�$�u/�.������F���E�	�,�MVt���NM�2�(�7�_��v���/� ��Un:���{�u%JҔͣ��� Vo2H��t�v���r�%������Gwn����7�|�Ƽ��Z����+h8�zͽ����`7(ks�sN:���WJ�-
�&B�����>x����D-�Zp4��ć��Ϊ<l�� v�����@åhgMod|��>�{)�����k�?dt]��ƺ`�s���T��&vD/"�(��ڤi�/.}=�8WT>��yO�FR�n���'���o I�l�'�����x��GB�Si�9�W�.Ī"�O�z�@��F�a�sz � B��mzz�	�ʭ��̗�j����{�aỠ|���StzZW�C$85�(�Jq�o$��g歓�n��Q*U��:~���iNŐ�J����Ӈ��'_H���@]�Ϩ�2!$�������^_�ކ��,�|�T�E����2�W�����#��f��hū?qtZʰ֥2��cŉ������x��Ea�'�[{���_�#C*%�3��0W_�X��l�z���F�pL�X·�%�����OC�����+C�+���A+�o���S	k�A����s��E�M:�����G�%\�v9:���.�Z��(<(��h��@!nD�6!�>�!���v9�K%/�n�o�ud���\QNGW �bs��F�i��7 ��O��S<��s��"���J��l���e;�/�d�}RU��}[�t�2��>P$D�����:�L��o�������c�LA%䫉���^������3X���'"{� ���B�+`h����Y��}�ݓ~k͝��i������u��`Wc��О,P�P��_�h�>+�-W��e�$��k��U��ol�&RE����������Un��Rb���$��u��5mR�3l�4�flÅDW���I�6�L����&F&R����l�#?���E�����8�J�Z��f���Fe��T����Dg&�y�Y���:%v�IWF��b8UI�ۗ�(�
������}�ng��r��*\�D�|���#
�=zzq7�g[�ǽ�=ݺE�\cj[Nο�a��eJdO��x�}*��-+k��[İb��3	�лNp��71�b�B
����_و7V��J���\�\T�Ma��sD
��	pej��=Mt��:�czA_5��߫�ފl*��GB�f���ᚹiD#t5oCz%U���3�68��"i�u9'D䉄-�f3QxQ�=˓3X�:����p�P�}B`��w��k���x�]=
_ݸ*N�����yah�ha�!7y� ���$��ۣ�v��o��a�ϖ��^j
�c����O=*�z'G���?^K�	���C�rs���@{�`��X�)�J��Ng��+S�̶���v�b';�f^�`�?sF��̈��u��5s��V��T,�V����?�1L��E������|W�W�����E���s�����᤟̖nӥ�A�*�=��/���dڟ�ҵ��Ƨ�y�=3��#�8���\bRZ�h���8E����������kM����7~a�q���k���B�����B���5�� )����>S,��[۪i��� �f�q�b����x��*i��C�8+0�k������L����=�m,�{.G8����L��nv��\><]~��v������]ڱno�J]���P��Ο��3�����1d�~��b�	"�Cs���*�1	<�z�/�ݨ���sl�g��\�����j^5	<�Rx�������ɋ�5L<��xc<�E�⍐�-��1Hl�7.R�{�y�м�m��^���Cņ���m'�o^n{���מ�$)Az�����
2�/-ǰ�������,dܰ$STC��- �i�@ٿ:�UnS��A9�s��F̝��q�cAm���nM0�(X��g�+m�b���r5,H��ّWq��ѣ�d�05���~��XCȠ�)��C����
�&෗�ٚ�ojޖ�M������8���F`ښ]�+X֢�ǧ�A#?ʲ&^Ȝ~��uP���N1����YԷk��J
��4�PI�:�G������L�q�B0`Hh|�љ(�^�x߂ZrY����6��~�l����]k=z;p2sn��������I�eS���7$4��ɤ3����B`Or>u�<!g���3i�k=�O����i]��j)�zi�Ĵ�L4�6΂,�GoT���")1V�Y5FT��먚Sp�>]L�?������A2(9C�@��Xk���I4k��t��+����]lnFc8�^���]���*�Vs�?�ɻR�t��'�Gs礫;˃��:@�_Y~Ł�T2��*{t�+�BIAe����a����Z��U�Q3�ot�9Y��/e�HӓJ�0N^�Z݇���\Y^Π�j�r��fh�#B���*��h�T���n�<�O�}�5,����C �)�M�'�:��k�s0DN���F��+ĸ�jm�
,6�9	�����ƙD��t�<K���~�S�3�}�h��Ā7�L�0t�r}��g���i�lU��
=�ݑ�����t�$�VC�v]�|@�2�o_��o,�I�~�P��HA�W�v}���L��-��X�\(jX@S���(Y�*t�p7����<�Mud��� ��B�����Un�ۃ���8u��T�g�`�yc�?3��_8�ʐY@���������n/���[�Ύ|d��+��kW�����ܷ�>����$��R�i
��v�d�t7$/���3�P�__>�����({��P$�\ݹ�k�T@�c@!�٠7m����V� ������
/�&��\uqo[m� 婛��:�7m*���dď�ο+�!�O
_j��E��<T���8�cLO�`h2�!�I􄽧y�(yǟ�SF9��� ���2^����������  �����@v�\C�|,,�2�	��KN'�i�f	�π��S?�|��@�V�m AwPݥm	��]��o���U��סr�{K�K���=�ZeȷIDג��ќ�]���քI���&��z!	�ȍ��Lʐ���m_G&�@>���Pÿ�Π�1���o�9�/C�[%�U��S�<��q|V��~��8Ś	�����ΐ�5/�A�f�\^�qS��@5*�����tċ0X1TH�
�[=�Šڊ1FdŃVV ����`d����c�M����D3lb�
Z<2DL���<^�ie�������ɗ?����5�3�;#��٤���[2z�(fxsy�X.��ο�RQ=ǫ(��Te��-�9�q�V8F��Bݕ�L�7G�=���L?��7�&lx��&�:��.�W�+����)�Nx�$���09L9��U��݃���	��X�W�>"/&J�"6���&�VW� a��nXH�CrW:q�KcR�Ry��I��wF8��?�u��`MU�l=Q�p�L��i'�h$��⊤k��|h~s��="df-��<E=��t���t�" ��E����7�|d^�����@3��e}���E}����rx�G��˲iX�ɭ�}T�Bb]H/�px�N�_�Hb��a��؅���J�������4���X���i�-8߬e�e@
v�[��\��ti�4�雼B���k����N�67\�ͮ%���桔:E�V�/9i�����������T���q��U�Q3c֯O�u��Ӏ"��蛶u?Tci��p*�%h�\N�$gw@+$Hډ q�)���=�TF��k
���@�@����`c�5�q^c�_��f(b6��';��h訽�D��/=0�����xi8fKhh⼋���vb�CEe�	)�q/t�`0娚jp'���Tm%��T*����[��(�q���'7~�)	\`V��U�ݏ�9�\�39428��c8��7�I�G��M	(�r�6���v��x��Й
�Q�l��q��[�Ա��`���7z6/P��cEaM�@SQ!,�y�CR���p��I���U��sT�B�}�S/���Х7�߭�!�෪����a��WC
XɅm`&託��؃V3VD��� ���S\�r�Uޯ�s��kD�Lf+߷X/�����(���=}��
sLC����bz��~�Af���l@w���&ˊ�r4��ҧ���p�7�l�E��P~ں����~%�d�*�͙Ŷ7�r\���q�HD���_����wiw^�*cR�R�~�;���^��#k�a��[��`�b��Q�&�T�f��׳E�j��bSꃰ�i/Q��vu�I.� [O7�Kk�/I�����E���G�1������QǜhC����^�>����F
�k�`ٯ���
]����Z���l~=Ô:v�ǁ�� 2�M� ����Q���4��偨4tt*��àߊا~��hw!�U�L�^j��Udf(�/ƛ�kx��!���
�[��3uy��Y˙�oz�EGz*&�ʐJ���L]�F I�=�|-~XMxT�(�b��
W��h���|51��-Ť�N�5h���d�pݠ�����L��rq,�S���T<�' J�C����EkR��&�Z93f��yH� ���
�D5��o 8*����EN�0K|�R(d�T�.0d������Ӌ�S�D	��ZK��ދ�}�*�9h���B���ku*��T���J�(�*�ӕ��X��+ �bP�^]"c�Bqҹ�"�$F��n�������^CDU��R5Qr�<s�95=�� ���D�ԇ&�$u���e�j�@�c��{A�R1�_���l�
����4	~ֹc[��ík�&8�Ø��T���SBP�ND��� �x@c
u?ʧ�;��eŕy4�)!$�N pa�ǽ���+�;���Y4�AҞ�{Y[Ha�К�=�n6h�A|K��bzp�\C����'�)�8��i��@�	�bFqr�X����=���{)TM���@;���ņ�O�w��=r�ML�teϮ*{�-�߾(�Xk�HTn����(�$A�SRk��4GZS�\2����,~8&�{�n9�~V�uͥ:x��zR PE�d?mE���$&f,��7��e��3U<�SlN$�x��%4��<���.2���Ν��HG>�DU��m�k�~�.����6˧�i��TWv��5�<�q6iC$s���t��T�!W&�f���_�ᐑ�_�=�����:I��Y�K�sp�̣.ny0Т�hx|��L��<'쮢�b�:bIW�{���o��O�.��+n'Ԡ�=#��p!ǒg q��myx�Q�)ٿf.[>^H?J��ޅ�+⮉�������w�T��gp^�b��g�m���ϣ�*s� 5��l��������7o6&P�2�q%�!G[j���,0�g�\��4����5(ra"���CC��K4�g�Ȩ�W�_��^��r�WՇ/��wC�^���J�ZC�1��N�F<�+&����&$�]��A�������xbEux�s�"��9��V��[z1������@�b.<�酹������bJ��W�F��_4A�~Vb)z��ʒ�.$g�n5�8'C�2O�ZHM�����ï2�>6;O(ͭ�D�a6ܠ͡�Y]�%K7�m6D)}O6���Q���g�tl�W��W��dX�1��ތ��\�bUR��ćV�8�����@}����I9&?G�Fz�6'������5��˶n�]��h�+~�
�"&��[�TɾjD�9���XO~
]�A�/���#g��B�GEag�7�L��o;��L��.�!�e�B޶2SZ�4�Cb��e4U~E%GH�����dy.����o���Pc�$�Y����{4��
�?������Q/Ӧ,��HҲ=7�HJЎ��ψ���#��Oe_L�J�B�0r��3:oI$�'��_M4�0����`I��d�V����[�H��ghL���
����=y��8<�`��/�	.G�����r7r���<1k�ޡ�.�J��T<s�K����RT�`�^Ϗ�OB�T�B���n��GU��#�������fx5��Ӈ0��xo�I!2�묽��v����SG��i�ˣ�Ms�=i�Ru����V��k}��XQ�Ax\.��Ւ����,�)�0�l�%S��G��w�`�ھ�U�
��w~�r.�P�^zۗ�]f�Һ���JbV��C�3���$��0<��z)��946����!��w	~x6�,s����G}'t;�
�]z'�<��*PU�hp�% �\A�X|����X[�PO���E��x���j!T&oWF����3m�+[�~�C��?t��tX� ��Q~Q��+)�U,�z�m֏T�Z����ݗ�a(�����X��idD�:ܳ�\$��j��Rr1�g�j���=���FbA�w��iR�#�F�U�8n���6j��[;¤�V�ZZ��iv �o�"F�I:RF�.���D�D�^O��H���Ξ0�U�lѮdn�)H�sN�*����^���R%��|��E���Ix?U텿kg,'�L�L_%��;xWU��e�8*��y����n���$����yHM`�!�,,�r�o����EC���Q���b�w�k��	j�{uϣ8��1&��u�44ߊ����/ӫF��h�ꡁ��1�z�N%�Ԗ{�wܖ.4�/�x9�-�T�II0p⠆����3���N_���
N�s4��Ѡ�r�el��c���)'85,��H�85�t���z�1HIW�.��`���3���"E/�E�k���{Yo>����m;(U�G{?/V��qv��-���Qe����g2�&R}V�\Ś�kxN�L��=�nNV�Зf1�MJ��
 ��ZLEL&��e���Q"l��@F·�%�D�xwM��{��_�> ~��A��'��pDb�[Μ��/H�6�Nv�VZ|�*��9�Aon��Y��|ʇt���淑��9N�3����7d�㬘`��������d#h���+�F��"���lQ��~�F��;���jd�*�������[�>W�l����;F��ω���Y)xz��2j�������O�~�1u��� ���}�X��d�H�c?;��Kg�M�}u� +��9��S5+�S���?��6�Y1�@+NR�)�k���h$L͎�4�Q����$��y�聜�D�m#�-Nc����ˤ���u�߅|�[=�>����R:X�CEd6Կa�t֙�����\k��?p�ڬ��8�pByX�#"�q�y��Id���k�g�����u��xг���n}Q��6Re@� h�hEncȒ�2U�&���B�Y��-�Ah-�H���P�LM�����P���_х�/�z����;�4k\�)e9#��׮R����4n8���L�/+�s/g�ϋx{KNA�#��b��È��7�qLP�>���4S@z�3F-�to�H׃��F���D�yI��z,әc��e2���JvH���ƿ*Ji�f�F�9씗���Qi�|?���%�u����Z*K��0�&�위�^4	x�?@�R��:��Y�nKM�z�sh�Mkt~� D^#�-���>Jց[=sLXv �W�S�X��O0����$>~*�\�cG��n#��9�a�:.�v���l�Ģ�?�U��(v�J.%�l'����8X{C��l2����(Jz��]?ܜs2~�G�ӠĻo$���k�\�9��>�#���(�%F�`ZG��-�+r���&
��,��]/����#�q�������8���j����f���	AO�����t�r�Z�d$Y�����\[JT$�����6W���?�ܡ�+%%i\��j�D���]XY������פ��+}����(@��E�zA�\Ţ:i�V��~�X�>�"wco�^=�{�p���q�NEv��;���C��l�IQ�\�!h���w�r�Ͼfс?ІtȆA	?�#�y�`����/uҦ�ˈ������H=j��co����Vڧ�*s���dēZL��UO�lHY:U���B�[�[��U�o@ֲxP�(����<�3n:Yu5�\r�tOŇ��0��a�=0/��Ү������O�93P���aР%E�h#lm�ȑ�|s�MwWǝ�R_��^�1Y���������ĭ�NsC���{��@�.���-����5M�	�<6FL�F	i5��Q>����Tm���G�t~�(/�^~��7A6����g(��"S�2��:iU�΋XM���[�Js��[��/K��D���^f�Ԩ(�>X�2��+A��P��e|��Ւ�@���a���m	z��[8J��@R$����m84L�%�PZҴ�H��򇿤�&Z+j���i��rzI�Ħ�_�;�����NUQh�}�����GZ�1��2�N�����@ x��&���p�&?�kL.+�8@��K����8�ٛCT�LP{�������Z��L��ğM��l�q���PP�-�������R�=1�F2�$ޡ�y����1�!(��j�l�%��㿊�Qv��v�BfQ9�:�OLuj�m��n�9��Ǘ�	ڬ�~���ku4��V���a��u���M�y!���a,[��U:�P\��</.`A
3������r�S`"Zx\�u�Pι/���$�n�L;.F%�ԭ��<�SPJ :��TD� �� 7B�Ә-�Ͼ��y�^�:x���o��d�qE@z;��k�Q9j^�.%ݖ{�e���J������<��n���l�ѕ9s�JYʒL{g]I)�rm�'
��OX�Jd���;�r�3IM�0m_���D�sJ��Uؐ��� b��6<TL�maj�B8`��E�O�4x7xڮ��r�]=G�Ĝ�<�T�w�Z�$ҺlJ�_��oL�����so!3R�M ��	/�EيÌ�1�a糚�,�N���Q���b�0m��)�`6h0f�$x�D�:����<���b?���	1r�����i1�]?P�c~;�Dܓ)���sdH��`�K��v{e�A��bUs70�wa�to��q��&@�؉�W��IU}�moI��D��)���'g�2ȧ�"r�������Oɘy}Dt�+>���Q�"�ScKZS�~!��A@���i����k�!�e[yӟ(1���K�P+�w5��������?
�@�Q�g�uw^9y�����H3ߖ� ��H�@�p83;(�L�6�[G�R�;�yB�b�}^A�Z���܉z|�Z�����-}��(������,%��$��8�}��_9nIB�S �`��v1�7[�AlX�&\�xJ�S>�����#�9$}⃿�vU7;h��#�(ђF+c%'��>KI*ьOMuU���	�[#�q|�`��'�&J��ԅAC-'��LI1�b��N��yE��Cl�'��l��#,m�e�K��\{=�q�`:
./�������B�;W��]k��r�.^nQ(���tk�mK���r�:S�sk����g�'�Z�<V��3����d�_ڄ��~ظ;!�5ep�X	^�ԫ���pLh!k'�jtOCa� C���wW��]W	=s�Ol��;��v}��blJ\{�i<���f��?^���2o���2ݭ ǟ�tZ��)�X�ԑܓ�$b�sm���]�bt7��H��){T2.�A�K�a<z�a�	����0;�2�m���K�-զ}m[��0��i��ϯ�(��B���ۋd��{sW�h����x�@aqi��vT�wD(��mY�]���	@��D�r��U��n3+�%����M\�s^����4G��ؚl#�}7��&p��s��u�j��y��E�!�:Q�{\�])����֤@Ɉ�׮�����D�m'�>x�[����;n2f$�%)�΃ |���s~⃘�:���5��K�J��v������	v�)�M�!��ֱS�_�xT6�{���ii���`b��}~�\��&Xbn4�M��F�;r3�����*L��c\/��*f��\+��"�2�dn�m7w��7Az#'w���|g{�7h��A���d�{�2�TZ�qZm��$L"15ū��K�ȐAE�+�҂��?��Τ���>���q?���n�l�+���Rue�O�����0�����Pg�Ɓ���/�-u>����>F�a	z�i��v�T2j�ڴ7�֡��� �ZLR��|l#����m+�":�n�g�o�0ʓI�bi�Yb�͑#o�C橯���a�]Z�elGq��Q�����b�)SEyσ���U�#���y��VT�/0R/Ҙ���o�����Jn�}B�UՓi�T����_n�?{�����P��=jT��p?r-.�o�X��A�F�&�N���[�V�f��p:ȸz�R��I�C-Ǚ�(����ܩbH_^sޔ"S���,R��G��,��	���g�;ҙ�b:�����$?+�ɥ�%�c��&F�6���Q0���@'��,ᳪ:mS�e�̣�&|��y�Jcn����,x;�3�֏�{�`w����ml�:�.��f��t�N.�f��=9
����z�[[��t�y�IRHJ��?;�Y�~����ckޚٸ��b���}�v��� ����y�B��!Ao�e��}l��@���)b\���1X
8S���7$��F��W���u(�8�&y�Gg�S�p3]�m�*�K%��{o]X`}����.��%���R��N�9�m>��������ܶ��1'i�H���S��wyޞ�9��#،j6gȂ��`0T4_����"�])!&��5�6��g(�Ȼ���K�_�޺��ƕ��\���x�t�Yp輔3����?w|��-���%�[����q�j�=&�K]h�Zk���{AbC	��?������5,x\��ֆE��/E=W�pz�	s���j�����R�`%�8�{.�S��+�75PwM~:ѵ�:Q��U�S�K�<!�>J�]�N����GcmuU�~jٔl�<h�+T�x����K�A��k��d;m����*�G��D�"��g>��w��D�I���U�YkL�� l�W�-MG�D���A(�T� wEu�맻���K���5����'�z�q�V�v��00ZA��PY������nE�-x�g-�&�{�'�O/�*: e7.����L��U�ts?��sɶfH2�b���!��H3������}��V�<���!��ݢ�l�5�
��R�6�&�O�Gx�5�[yB��2A��)�"���"Z�pܞ�h^��I�A<y�)���
_)�� ��C>ՖOo�x�<�7w�Y`�0}�H�S����!�S���.6���5拒D��'�3G���n�5n���ю�C��@�Cߧo���ϩ��'>@rKQ+�|�R�z{��H�m�9 ܰ������kK�����++]���O�k$NZ�l��O(6%���.��6dS�i)���ss�wR6Y�HCt�0Ƴ��5��b�Μ[�MSC��V^ُv֘]c��N�pJ�[E�� ��-A��A�9<�j���Gq����|y�,���<i���V|�޿0�_����n�V@ 	���!��VL�����M�*�p?��نe�x��;-��:�4Ǡ#�R����"��!upM6՛=5pvJP��F�cn��|ڷ@c�\S�8Bd�I�1b?t�<'��|u�2=G��Y�l߅�����oى�w�^���؊�|�E�ѯ�{]]�^���� ���~s���F���cK�f�*�	�������r-��AltG��B=��-��$ѷ��:������q-����}�Y�����~�8����r0��yF�/GoVQo�����Y�S�=��Ձ�h����.JYE#�H)ls_C66�?9:G�Z�͍kE��D��nQnY��-jC�(�4��,���a�����o|dX���Όh/+�`o�lH�p�sp�G�[������т�P5�x-t a��\}���䦔#����s�OR4�E$5v͛d-��>l{��Z��?K��P��R�o�C4�ʹ��VQ��}�ug���.fV�e���^o},�u(G�߅~$)�A B�;X��J������������Ы����t��WSQ��:�c��� �'x�|��E>$y��I�p��$d\>��3fkj��~�j��{����T�����a�BY]���>W�$�oT��/|o=��'��XNd���(	�]�߸�oĻ�͑L�/������U?�B7`-�V�<�E�h�s���)���2k���A�4�P���r�
&��#}�40T����~1d'u��[�tI(4=��T�o6l
�d.D�Q��Z����
׹�{ܺp<h�)�,��6Sz�֗8&G�IIՊ�cU��W��Vi_D��?�P0o��o�uVӺ�S�ȏ����/����R�v_���9���
�R(jDA�z����/����C����6�)T���O �����Tn �]䓏�U�9G�<����>���v���f�Í]y B�/�B:��*G�E��ע^?����	���R��� ��[k���'W �ǆ���΁����M�_�
�;;�/�l*'٭�� ����*�,�/���A������F޺�Y�n�7a��>����·D�A���'�����RX.(��
�c���)L�]��Rp�-�W�t����(8?�/(�"��5���N4����G'�o�icZ'pd��JҼ!^�M.3� �=�D����ͳ�'Kb��+ȠQil�yS9w(��)|('���Q���>F��h�(��$���Ӹ��7�Cۿ I���`-@C+��x�MB�J*wzB�0E{�W7Pr�I�� I������^߉t��cF�	a�{�~��M[��p�b�