��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&��n?��1ů��> K�-� �&�T�Ek/ֆ�\�놭5�DꢘP���+L+X�4��J��#�0�8���������l��jT��+�(���������6�MC!D�;�m�퓊D@v_p��䙋ⲝ��C_�6�Ռ��#�� ���	RD�4D��畓7���vn�H���0���fX����4 �CS�C`{��;�L����li��� y+����FD�p"��]���y��R��K�({� .؜M�������	^5���ɋ��&���&�@*���
e�� �t+���
_6��O<��7f�M��u���m(MrN����z�jL���@T`��M3��c�uQ�Y���%�dD���,�~^���y@Ga��(����C����	��G�86�S$��ɳT�ز8���:r��/y�[ݦڍ#A�����i�&<nU��<[5)�Z�-Ĭv���0t���d���"_���:�'-��d��*��q����_d�y�N-��~";#��������Y��؆���	6ZJnԷW��έ$Y�K�?�4���L�w�Wmiɶ��Y�?jx#*�i���F�m�E����O6T>]i�_�9;�!(��kH7�OS��_��[-M�((��lO�s�$�g�x7`��ZV�E���F��,9�j	@���]}<�ahb5~ãdl&I^�	v����-�@�@���	��!��d��`j[Q��� r��;f�i�.�m+UH7��/OV��c��������l��i��M��*'��?���G� SK�M��H?�ç��q;��)��Rȩ�"@���r��Ml>8!�S��L��EgeH]�8��>]GR=&���C��i�Za�z�,�F��h�q��^���wT�a���%�9�n��?~SИſ~�mu�OlIv�4'sT���/a��^��9��*��G�Fh�DM�_��CN�<�_Pg��O5��}s�%��m�o߫R���X�Q?��dK�Z|:�=��y�P�)�㿶$�6���,���S�E����Y�.*_P͵U�Q
)�ړ��N<H�h�F�UO�M��V^r�*L�3獝 Y9C�'����ҠbW��̑,p_�Hi�i�rU�u�"�-�a�9.�f�'�fct9w��0.Ht}>`�NN����r�(�f\XE}(y�;��|[�u��ߥ�\�MIu�*��@��Ԗ�?n�F6��&� =2Hhg��`Z���E~��	��DH��7�Y��7�:Z9��'l���AL;��k��Ȇ���C���Лʉy\�$[Q����6�͙A���Xt��>¬W�:. �#Y"��{��?�l�i�_�Xӑ�_lG���F��[�ҟE����S^b�!��Dy�*���&|�g��^�"�R@��~�IL_]�#���]��{ݙ|��Ax�Ml��R-�8Lf�V����>����ưi��G�+:�OU�+�y����6p����%�f�!���^6�B�	���J^�S,!���%��s+έ�;�4�
�7vd[�xo����Õl�|�&��r@����O\��pL`���½�2����3�[�x��H�1��F�ȵ'm� T�c�뭾F�wVJV�XI��p��j����/�",Dd���^6��L�\�O4��Β�\ܯ\6&����
�� �.,"���}f��90;.@�LZ~0��O7k����7w\����,L��u㨨Ϳa�sq6c� �*k�H�(T]~���]��������MJ�u:�o�D5�#�#[F�f^;AMMq1k�CC�G�_JD��"���E�(��ش{B��Q�[�?����_l���n��Ù`���L�لA�n,·���V��]������aԍT�h��;�/m��	<����7�3�[_��uFC���Cb���Ữ&@��B]��?��4���S�$�_)Q���"6���e��E�j�fO�?KL}ln<��k�nS��4� ���* *�(� ��v��/��hW�~�6��u{Yl�+ج �!Y�a��KLF,q�����h�� ãJ����-�[��l9J����x����hXo/}׭�ؔ�M$�k�t$�i�hb���T���l8$BCa[|��	�m����CD)%0��X��<�Bs�����������]m�=-�"���i��PPs3���t8Y!�h���b���\��e���|V���iOCT15\�e#6haVЍ�9H������,F� �VH�����&���,�w��Ny�̤^�%��!*~R��Y�^>W9�z��$(�\>=�$�O�������SP��A��M����A���n�dzi���Y%�Gvc��c'Kl�=5�Q�:��ċ7��3fb7.!��^h��_���숖ù��
��ʺ\P%��6�>���9t-�2����6_�ļ���
IA�>)0e��E���ݦ��������5����lX|>N�(�a��ǴH��I>������J9���^��ħ�P��_gGC��3�������9y�ް�y3�Q��r�T��8�jǜ�o&�!O��v֌\�ev%+��K�JC�&l����� �sd�uOg����Y�m�}��]�Yy�qz�L(�*���B�՟������� 4�WA�k����П���?�~He�sΰ��v%�J�nҽ	����w�����.<�_���W��6���a��V���,b&|3��7�o��ZV�8��N��S����W	�S�A�vj�S�y�u�7<v�8�k�~Q1�h�dh��mD����M�$Y´.$�9>I���ta�iq�r������Fb�d�`Ѫ07�U��S����Eyg�`�=����\]	yn|�nL	RL�Y��FE�)>�w'�k@=�NG�[�#���Ʃ�6�����^[�ݏ�[U�} ��@`s�4"Ȩq�0�������@֌"@�&Xen���J���+��r_Ґ������^60µ�/k*VhA�����8��}�3A��N��������b	ZSŹ�hB*�"f�/ۮkQ��"��=
rp��αQ���\B�O��6�v6�����a�F�n�\&���sza�`���[�U�!�$߀����� �.�U]��������
�ᬌN߀~�b�_��#�.��E��Wd��s�� �-�����-�80)Uf������Xc����R��珞�Q�~6 �"��l���X�=��s��<?u�&�f����X �u�y��R�6�R�-sT��@���O�௯�:7�L��q<��P�i7��#E�j�a�׎������.�N���z6(��ΰH����:g-TJ1��@n��}Cj�t�����Y�Љw�KJ�ݛ�.�.���l��is�q���&�q����1R�R
x�֭u�Cǻ��ڈ����^�L��Z:b:�"xn��4Q�Ǯ�����{�ߛ�L�����~��(�W�ǃ0�G,88������<��"�g0I�*����`���/��B��ڄ68�d�X6Wt�`�d�٧�iy5���]�2���U������`w��c��U����p�����$��"_����8���i~�7�v���]��5�SF�ʿn�� �h��RC��gR�v������0N>�ڈo��{�:J����j��S%�֛6�_����*]	\��c]�{Ý>����ANɹǫ�.we�0��Y��%�%�F0D�-�l�l��HF{Be���J	��%+�?�
2-2M��eSFw�9��r����*A '�d���sY�U2ԷӼ�ڠH,5��{{e͋�L��O�6��R�&"md�5m<�	W�'���
����B���鯦���5��4B�j #�����'��p�aS��u��-xQ�����Z�k���@?�)��@��Q`F����2�J���x�>0eK
[QrϠw��" 4�ȇ%�F���ņ��i�7&��)���K�x��X�[-��%�U��V�������8�KP��D����u"��(Y��B�[37&c��[���F���Ńl��� �Ȏ�s~i�(��x�`_P$�}s$��h`j111�^��0�6�8݌�F`�v�����8Tj���[%��;����C%H�s@��7d��o|���z�ė��%b�L�d3Tv�H
c|�*��Z�k��8g�bŲk跗Ta�59|�nk��'iq������#�?������*��W�;�Asf�GuBa��G*~n���/�ܠ�bO���3�0\�~V�c�ñ�2�l([B�PmѰj*␪y|I>m,{ԭ�Q^��e���ؐiF�YA�j�I�	ѿ���}���a6P��cd~��l���1����fx\*D���rG�{%���~����":��	'\�⸌ �1�����+�+,�S-!���< �@�-z^w��|�TZs�;,ٝT1��]��Р��#���
0cD��v�s��s�F���Qld���\
)N�����u�4�5v��\�����h��@���2H �܅��#�쏍�rc�/�K��u4�H�e6�W���GJ�QA�S@��୫�@.C�q�A�a���,Y��X�,x���EI�$	�(�"�L��g�Cc�9`�^�x�!߱�;|c{*��R���4�����]�ψ���C��u̷��ޏ���C��B�DG-X=g�}W�o�p��+�@�K{�J����nֻ��u���M�U�_ov�;4�}��:v��b3d�0	��Dv3r|7ѵ��V��Ny��t����T.x_�2���΄��v	���N9�Q��J@E��ͅ/��Z��17jVPR�<�er}X6R� ;o�^O楂"G��387_�K'�N�j�+3� �Y @6LS�)�d�<Xj��Ӝ<�k�P���8�Xa>�+d9�na�90o�f$F������{�^�uU Z���$�}�xgez%L�^<Y�OC��]e���M��p'�\�EMX.������{��2�Su�S��` �~e1�������X�\�n����{�%����v� ZMO��O��r�v:ɣ��b����U�R�um����Y*�Ώk9Ih�PN��<�;�s"���F��f�ˉ%�X�n|��Msa�����H陋p0�4��\��r�� 
%�������,�쨰#�Gj�{�v��:IP*B����B	zh{m�)�Y�KA���z��n�5�^SN�	�q����_�rig�pBH�P�(j�mDH��]3�������x1lvu����*S��(�����g��P�s�Exv�ov8�{�ܘ��BgZ�K��M�O��<�摈�ڏ��Z
��d�����o��:Z��o"�*�
Eء4Z����}3r�xw��]g�Q��H�b��J�# ʈ<#�����uE���wT�A;] o��7��h�0b���4a���E��r�d�ܿ��(AՉ�aYr])��ۍ�H��GT�}�d�&�C�lT��Hh�9E˜��Z'����Ϻ�o����mDrH���a���bmAB��F6*��d����L����چ���9:�z��.�ų��[Y1�/$L�*�|+���������|������\b�Y=2������R����Z��:��Ҁ��6�,���7p�Za����~�(+�pE2�i,��%�R�;�,Bȣ
����.�u�$�v��7�"����Cg����LD�dE��E}�Mc��T�$����`5Z��{��������{�'y��=U�A�b����^�C_vАq��)�;$�tb
�Zu���?��e��W��&�Dx����n�р��+W��.�{��u 2|����k ��:���D�eV#��9Y��ȫ��t�Q�z�\�xf�ߠud����YW�,t�|k����V?�I�W(�$`����n�2�����,���s1���} �$�v�7�f��Z��r��F+�k�2�d���H�J�ni�a���]@��d>���
�V|<�x
U���q������M�^C��W�h��q<@�e/^�'�ۦX�םyaJ�ނ��,��%6����wDVh_�JF'��jaw^�I��bmQ�˯����с��&?�P�A�FP^�ȥ�M�P��L���~q���B�_ܥ	;cz�)j��le�H��|���~A��`��w�B9��������-�@�d����e�g�0ɻ�h���5��)4v��6�?�nz5p��o]��C%��<���o��"b�Ͱ+����MP�0q��u��w�ټC�a���d��5d$� �%�]����UImW����]�_vK�:�D�S7�r�{|g���0�M&�7��k<�0�f^&	�k��̴�;k_�&�r�R� \��?��!�">P���k8l�����]:�o��&_�<�̓�P��آB"�	�T���/�-��KJ�NY������W��+?��Js����Q=�AŞ尖���� �(j���oT&��D԰
�����=+mN|���#�K��e�*�D^и@��^�r`e;R5K~"PCR�2�j��\�<n@m'����-a�X�:B��V�kN�@c#%��r�oq�<���>ʗ	}�����%s_�!�z�EH����P�'[�=F�"4Ǧ�0Ji�.�4Ix���}#"G�PV�z���݇���L�����6�0���m�mL�u�����믦���V���[n?�>���!����ݔ�� ��_����(��V^<8�>;������T�`���v�T֓@�>Ǝ�n��񑴧��h�K���-=_grU����c(������Z�RФ��E�\�}J�����;A�ou���.��(%�2|�Ц�7ǀ�aw�������]���k��D/
��2���6_#��I�Й��L�.�#'��H�V+d�O��FJ��9N��yb���-h�������1�)�2 �	9���)�Z�T�j}T8Z�t��*0j@xҦ>�q��ǐ�(֫��o��jŖ���A|�����ޠ�X�չ�s�Ub�� z���P�����F�y� Kʥ)ٗ��#G2������nu>2�)Y"��"lI]�uG�:�{�3���^=8�[Dh`#Y�`B>�Jn�������X� �[(H?a`E����������ޯ�Z�Q�w�~T��\$�%���z���Hb�H^��Lu��q����	F��Ou�3�E�U�Ό�)�PA��Z���k4ؑ`%߻?d1�O�qz����/�����q��X�_��֫hKd	��F��L_��)�����C�u?yWג!o��!�dR�o��h8�`0�|߀翲��X��uC`��`3�/��؊�*S���z��q'�3��{1_��;Qη2k�,�TIS�?@P�@����C6p��)9J׋dN��%���r�W�/0�6�I��9�F���Ә��W�i�R�e�ijDs�.f�gp�\��χՖ��[ƴ�T���pJd�ϩNZHE�x��[Əܮ*���1
�vT�!Q��?m��1[���C�QRѣ�8�����I�0ò���ĬwV�����ޮ)3������� R�ǉ']G����.枤^ǥ^(�)�4��pDY�WM�|��z(�������j�&��F�U��D�&R�yy��[��#��YI�҉��w� �����{Q��4Y)�I�o�{��W�9�(�%�E�e�5�A>������ToX�Mia��E/Z����'�6�;,�li4Þ}t���k')F���J�O����"|I"Z}�xn����G���.���=Z{���r��U�/���J�`�U��S�r�����K�͂,�Xd�(P�_Q��]C�����F �#{�_Q٩N*a�z��[��(�N�I�q�N�ʪ�T^j ��������r�D��:�>��q�1�8\$�,���j� 4dѼͨ��p�}ֈ3E��v_~�n�Eζ@#{���c3�>j�A��������d�<��mR��mc�lh���V������꾂 �̹���j���g6֬dΞd�b�&x�IFk�"F�4�ڇҰ��S���c���7Ⱥ�T=��&Uu+�Y����N�΢(Mi0H
��֫f �'�	dNy�{��2�0Ŧ���^Ӧq�}���D��&+/��p#�B��#� _��u��>�T�(��G����Ti��^]H��v���h���An�XБ���0\��j��Y���(�fn;ݸ�m�-Jk�ֳKA=
����B4��o&�x� �Y�e�%!��Ui�8d��o	�{��q���*&f3=�<m��K'�ѫ�#U��F�=�c�5�̯�d����V}GY㼁QƢpq���Pubj�'!�>�Tk���HT#�9?(����0�[�y0���Y������̣1� -mϔ�Ϛ8���Ebi��Z�)	y�b@�
�8Y��{�B��Es������'ϵpS����({62O�Ćii��G�p��$�)��- 	D�Gc����bŎ������16������W�I+�[�K޺t�o� ��\�-�*X�� �6�}�j�ax�T�.�ϒ�qi���=�
8���������/2�#A���L����p���-�$�{�G��V%�"��iYm;��jk��54�/��tH�6w�q���QW��
΁ 2�Z�(�~� �o�����^��WjХ]?iqT%UהO|���p���щ����*U�ʬJ?\B̧�ms�Tj�]�wjV ��N���	}��$-l<f<�>�|ƞ��o�uJ}��gs\��1�W��Ô��7��4h��4��Uvw��d�j��{�^�RV��G�,���s*t��@$��/�d2�w5���JP�ȖzF�Τ�%x,goXrY�˪4��Ѽ���ћ���sك(��{`O)%�iD`<�6W�(Cniūt�9���(��4�"�G>��z`N�kֵ�o8984Vb�Z���U���W�.���ȡ�Rx��+�nQ�(o�ٵ���e�8���<;5��j*&�٠�|:�
ԡ��d*=�bc@`=8gDG�����;hm�_7�4�#��E�D��L$%!Q�P��hC��%�W�	nl!�����Na?t�	<�؂GxN�2i�DD�j�d��c�e[΢BC8�Wӓv���!�������1a8�K�"$Ho�ǟ���7EHF�痑pn<ߌx��?�h�)�U����L�z�P�սk��Y��L��l�����1���U�������FD����J�dW���z����WP��Rzط������� ?o��m_����jU߻�ӟ�#`&^f?�v��=�{,2 �[�q�Fmh�
�{�Z;l���J�!9 ��,���ZgҢو!-�K`=�B�3�N�ee��rΫ� k���ğ
G�p�2� �?	���/�2�L]�|�Ic�9�ٖ ���\߹q�-ϙs~U�*_��*�[���@����(X�?8�f��&� ����l)�����~����!C�PS��?~�]������4��ыo\b[���Pߟ���j�	�D�F�\�=bV��NQ���_���+��N��f0�+�砩�3��{Z�.�i}�ًFE�6xs���������>i�`j�}jE{4���3e�1C��+\w-�2��t$�T"*�R�!h\���F�k��A�KSy�� �����A�v�y�'��L���.=	Ń��+�Le׮V0��.���b��t�B\O���,E�	.����Qِ�Z��'w�2[
7�����G8o��thc��s��A(�b^�&x1��~,��3�/���<F;�l�2������C�9F_o�|ᴠ�F܋�`��|t�E������}ڦ�t�F%(�]����41�4n߉NI�Dݤ�6N*��i��J��xH��g
��"l���w'��
��� ~V~����{n�hk6��z%҇�f��O�ea�!���'�5=�s��X��#:��X
<_ս�S���t��wH��Ѻ�d1kW�ؔ�v�n��yE������'s�g8��rJՒw	�u��g�x�O;>��E�L�ף
h,�1��9�K*�С$跧� ق�*Ĵ]<��f3�wFo[��K�Gϕ���o���� �JpV��e������w�PoV�
󯪥�
Y�`oF?��N9)���Lr���j=&` ?xÒ6����x�g�w �R�0�Q��:��%��~[L��U>��|7��w星/S3ʏo�F����!q�7�Z��G߳���L߹Z��?��8#R��T�~{C=A��,\\��/�@�p갈Y�C���<�be�c�18������Ӕ����34�������8e��g��V~��m�I�j����xf�*��Kw.w��Î��u���hNQ[̓�i��S��P�B�� `5�3*���+9�g�;��~��/�O]�˳���!iY��b���՝>ԏ� �Hŷ��:�ҁ�/��z�K1�f[�pyjg�G��u�����D�⚂��|��Q�g�O�V� �ޖ8��M�}�k��(r�K��x�~�d������A�yCJO(`���&8�MM�ks��\i�{�������Ȱx�-�Gs~L��\]�r#iy�d���$��~Na���ޗ8;�&]qAk|�	ỷ�GC?� RE�gJo����-UR�tB�\����K4��ɫ�I巡������ŅI�[���@�l�f�أ�ܿh1@�gE�y�\�N��	N�@�{
�}�A$���>�q�'��f�1�BE�w�{1��$��K >������Ρ�ξwؗc�CG@A䉢-[>\CK4r��lM�SL�ɺ!-�u��Y�x� �7�I�sT!f=WY�䠜G��
0�X�~Ӻ�+۫�Tv�'��R�
@x����(#^��|f����dKWy� �C���e�7��5
��W�o���&��%V���t�At��.�-+٣b8C*���l�u/h��M��bK�S���~8�&��֭i�A���a%���.�p���k�
߾�w��}r^�s^���v�a�:���Vɮ$�۳uhCFmŤm<�D��Ъ̣:��S/��)â0J��.61Tp����l�����I-�.%��ش����
��>+����R��g�]lL<�\3��f�����ψ�5��'�p�g�FT�y~V~��j��,�o����}$� N_��&5�[��N[�h�O�����UAլc��gD��H_����ܳʆ#�˚~��1���^�Ǥ��oWn���O��޵�2�q�0�Ù�I�:QkpG��ރ�y����z��
fqu�:.7�-����i;o�2q���M����|H�x� -4��r�RF&���ŝ�/Pkv��!UK UΘeg�d��j*ȩ+cА�ā��Vb�l+)�>�)o�S Y%��f6�8�0�����Hj�3��N����5�Po���zK�H�K�siD���?�ܼ�G�{A���7
�o��|<�YGFR>�T�Z�}ޯDÄ��k�;]��A7�Zɏ�H,K^�0��#*{�"����ɉ�^�\Ҙ�3�n}�~d���Kp�Ԉb�Ѫk��e/�D�i�_ A=��)ΪZ�L�>�����>�o ����OZ�C#�Y�K�~���}p9i�}iL���}���J�<�M�v�k
��u���7.o��vF�d��a����t~���M��uܒ�8��q�ȉ��T�5������To�n�(/4��v��g����'%d��}�v�l�F�KH���ЃIA���djU��e���,s�J�i�7E��5aU�w��A_�2�R�Gɨv�h�0hB&˦��9b���o��+�0h�d�l��-n�����j�˿�/N5(�%T�ꇇx՛A��D�P�����y���ĥ�<m%��9�憛��L������j���k���w��N!��ט�WZ�4r}��Ht�=�x����Xz���T��W�P�D��U�OG�4`�i�ʬ��Y<j���� ,r�Z�M�!i����6��)5d��+:: th���{X΢���\"����i�f"��ф�j�p��ק��Fzv�˱s��7���a�'(�e��J7�%�F�ms� s�\
���%�_`d��=���>�pN��ҁu��Kv��)ݽt��N�٭v��7GCd�F�G7��i=zZd�(HNq��8�Q�6�D���|!�7E�>������{|Ϧ�9�Id� N��׎��)�"x�����������5����>�������2����4;=օ�=9���_��%T	N&�����AI��T%�ߌ{����5ʂ�#�R�5�X���tȹ�l	��R��R����H�ȳ��Z��^n����C�d��e�:<�a��J5~T��"i]��E5�5+dq%k�yx���ݽ~
*1��ΐ��~+:���:���J�D�ɓ��qV�
��{Lq���,���z_Vױ���%��2��f�i��ѽ�"t$^p=�"ѐN�h*0�#]�����m��mj��M	Y9�7�+H=���������Oz��VKk'���T����K_{u�[@�~���+��l��M/?�a�(���9��w�ݚ�RBNE��P��4��8��%�\�=w�d�J�Q��l�m��/d0AK��S��h��L̷�ct���h�N�$)�je_9��0Q�����ƹ�3��l��&�33��D��1�7`�Y���5�	?&�'��Z�V�4hZr,Y7s������aD���nH��q;���9h�0��g��~��N�W%P!�� �����Q|���[I_+#'�����(.b�d�/R����A�œ���Zj���am��_���W��Q|k�kk��2:G���J Yۇ��f+���O���W�o�q��W����l��l���}쨘<�>z6\^��֊��.����0�5b�,Cc�2q�$ �r��0�m��-�啤��������lDX?� 7��2���!BD�h��>�/����\^ȡ�FYn��������b?3��ѬA�.�c�?Os'�z+|$�-���U��Xcj����.�{n���6����ta��x�����kI�7��p �ޗ$�|�%�>7���
p���1�;�D��*���`UT��pw�ӯ>0{&�eF|l���瓊��2���悔�cϰ�t ��2�����rg��x��+��!N���x�c��?.��R�@i�9~���$�G�����}䁑@E��`�ݖ�b��3��n+�↬����>��?�������R ɽ����+q�����:v�֣v��B�!J�P@��:���Ϩ>�G)�;v{q�=��CZBW�$�&��3\�mE�M4�ὗ�T`s�ߑ*�9B��Ck���-"/+�� }D�5 IL�~�ȵ����-g�
H�M��u\�Zg2)����6�����\@�y�r�+˼>���p���>��2.r�:�\���HX�)i��Yxd4��-��V{WU���l�)�v�+��,��i�����W78�/��?�H��b�����t�=vNa�G;Td+7:T�;���v�*����'vI|&���\��q��ۖ�V`3��%K�pۜ��Нo�ֲ�9&'�%J����9az�K���܌�*���	�;�1�s�4J���A���[JJ���bݛ�+��%�f����f?�D�3��`�뼰c\�'��~Cg_ lߪ��J����C�V Lk�xsRA\e�u"|,#f�E}�!c��t���Q�T�ވ_���?x]��6��װ`�<��X��%����"�`�����[�LMQ��G��g��	���ڸ�3�b��H���
��U����6ɬY8�C���1���oy�t�v�8U�@[~�����zi$�&����A+j\����s.���v	��P�T�fq�|�����WD�ّ����砲"i�Z*�uS�S���۫���Ð��tB{b��e1ޱ��ӌT���Rn�*$�3��w�X"�F�t��G��}�
���|x5����(�\ϸZs�i���ZV3i탠=Ry����IK�r͓̈́�����NR1G�?'���b�y�R�I��EЬ�v��I���:!O_x�$��A���ф��_�}��/K�#+�����0�Q`Tq���A���3vY�s��g����R��lB�`�:��rA��=��Z,:s��V�moT)<���4T�`��H��M/G#�]�:z8a'�EYs��A^�B��H9��FV��M�̗D�Aq�.{����~��"���j d8$�oIf٨QZ,�/�8��n�3�ţ�� ^U#j�r��TL���}��hm*\?��c�n���PϦ�8��M�4��yb����s����N�P|��t/�ħ�={�j��x�9�6����D�
`�W���w��XB}�j��D
H��Z�`}����mCʢC�ZX&(?�6[�=�c�3�3(���%��	|q?ʝ���2%�5���4r�&\dMn9���ȢM��[�N�Qc�wrE�i�D��(U�}�	���7Ű2�|QO_�2@<*�.XQ�r��do����X/G�G�ؼ���>.�j�4%qP/��S�a1��r0ޚU�����$�E����3���� e�$I�G��ϳN���R��_tq�*�9�J6|�ˎ�"�?�(UW�.?�煥F1���[+��'z2�������%��z�i7�J:u)�J)����6��T{��6�*I7kF�|(��	��q��c^��;x٭f:-ͭ� �U�M<�9��m�<���E�}�(S-��אoBn5���LA��s3Qp�H]Oڼ���$�$���x�����碰��j ��@R���6�܅2	(����>�`��"*�e�]��0C|���4Yj��5R̀���A}�.�f�og�iy(f���g�nU��XZ~�>���`�'D�R��p
�����Ӊ�y&�x�w\�i� J����܎��#�fP���M�;�d�۸�_��-�~6�c#Z��]��Ū"T���>�DcY�^2o���������\�ݾ�{{�b9���!����8G��@�~S���P��6|ߣ���n(�n?ʹ*�*{͛����Fݔ��9�j-'l�Pn�7�˃p���Y�J����t�����k �mz�8����pR�]��3BuN�\�R3�
@IҚޝ�oz�HO�V�*�>o�Ӵ����A�4d�X�s

�8����?��8��O,��"����ӝ"��rM[ٴ�H�X��|+�{|]��j��g����N��P+�Lt��in�Tf��Oyߪ0z_/pE�kVwb�V6�l��c�?F�)z�F��$�W��I:�q$�s"*�\��(��7��;��B��F9VN�|�i�>�*���2������I���|�􊸣˭&���A/��&�(���
�P-`x��e�A�+��f�A�G_Oϻ:X���1���ܬ7t���\�\vm �C��ۄB1��#�+5�7�<܂P��O�f���k�B99�R��!t���v��/' B�6���/��V=㌌*`���2��|f��s��'B�=-b�ЧerA���(%��7^���5�VI�3�LU�pj�Y����-Y��\B�/z�~�<q�@8��'��bs�>? �MO��bH}u�8 (T�bST]^�O����q��+�޶!�(q]�9R׍�q��v~m�/º�V�%��T��WĺL*3���F��2�o]��f�)p����Of{���ef�f��K�1F ���B��|��t�w�*r��&O��������PN�=�����(&�����'c���"����e4�*kٺ�6)�,i3�A��>�5�i�zqH��~C��Տ3e��c#7%Dܖc�trQ�-Y�<.��n�v������p�guAAC�I�o^v,����ZOH��v�3��b�i�:h��B�Ǐ�)�X�d$ﭥyn���r�ws�7h��'>�6�f�}F����Z�Q��#�T o�K��+�<�Y��3B�+�3Lz�$��,�=�}�I�hI+@}X2_��(T��@�=�6M��۰tN,u�̃K�|>,����1�d�D1�B~���e��,�}�<�Kq�,�Ҩ�)��o��
L1;��pҭLk��ɷ�����N�iD�1k�;9ǧ8#�{��կ,��[I��͡C"�V��{�k@� ���Df֧����w�U����T�"#�>��H��k3l����f���APaVu&�r��Z��➥ ��4�z�G�T��]�g�Q@�q�*9�.a��x{�b�M�
����|U6�&�*�z�`�5_��T�� qבx< �7��Z9��쟕X�K/yB��������3ͣ;�HG���Uh�?�C��52
W�s�;؍b��Ok�]�ڷ��fJ���f��m�����0̑t�ZC�?��u%w!ǔ�t5C��yŭ����@$�i�6R�+��B�"����yi�2��4��p^5}
O�����T��ػtAsǴ���z�Ǯ�ӹ'����A�u� ����+I��j9���H���B �Ә�l����/��ϩ��8�ϏK�:���8}��d���eF1D�s���C���A��U=����+:�7�qZ��c��4�-�L�z����|�@�B8��2��)�Y_@D/ti�8ӕ�=�ָ�9a���(��Hؿ�`�t��H��Н]���7m��|��U#�-GS� .1o9CK�c����~s�H�K�¹�5�Ҁ���w?����ۙMdsϴ��dZm������`�l� ��kT��0���N�(���4�P������D��C�?k\�Z�
�4� m�����?�� ��A�r�q����Ϣ����2�qI煾HƟD��(��D��1������hx�O��	� ��_xs�7�]�ZPf�s]�\�Qe3�G²=&�P�A��3i��="��)�6�F��+��G��^�1g�H���H�ܬ�z+À
|E���Iz��/�XYbx�װ��6�b)S�3�5_�d+ѣ���p�N�1FTʚ�O�lN�����3 ����)ݹºZ�<o?E{'�{"Έ��Z��9�g� 9̴�{$�@��������+�Aķ��24�[oc�Z�B����Y����$T��������Rd��P.7'0t"��[�=�5�3+`��`�`�+�a��&���>0�ӌEQ�˽/���7������cf8i��Ҩ�(2�${C���p�hrIIG������S�r�Ɍ�eU*�� �j��}z�ԉ\~� f��A�%`[�Io����;� �aͭ]-_���|'���{�a�֛`���s/4�c�q	M��記�����n�V}ƉJ!���{ơT�9��l1!p��q��pstb#���/_�>���3.L.�\�i���uvF6��&����!��<�V�(O/$<�|�i�2�`������Lm�K؉�=f�e�������� �����ܭ���O0��U8Q.����?}�0������K{1H�GL��,���"�[v6�O������b��:}JL�@��i�)�\����&Pƃ�˴�D`m�-W&��'x;��qB-�f�v,��ЦT���r�+K���F���S���Z�Ѯ"z��H��eq�ь�A�2#Hu�)����?���r �U8D4���4Z�QS>��VC�|�j�V��'�9��7Z>�><5U�sD/B/�N����-�|n��Z�ڴ�tv��z0 .X���������i�pFHl����)RB���1bI;��V�D9�_��Tť�26���])΂��_J�M[)��"�ZC��{'3��Md-�����gt;�&&+��P<ï���(7A1��<C-.�aj�b��C��*���k#�Ȱ�?|��LT��k�,��	��C�?Z2	�,��n6W�5�q�������	}ޟ�8Yr�ٚ�|��������%��O��R�҇(nBj`�i�X�`j�����Dσ�5~�v���J��X�@���k=�U�8�9NH'=)���� {2����F&Ɇ�mh=}�g�o�����d��;DQ�WݑVc�mB�*9�p��zȮ%v�Ăh�1�߄�����@ճ���;=gH��U_cߎJ��5�Bq��@�%ғ*�˞s���apD��\��;�<�ͤ��8v��o���܍�,)~y�E�mck%�QH{�-(*��"�5_���������m�϶�Cuz��T�[�����<&����<d�3L	�P��o6Ǉ=򓔘p9���f=4������;��,�
,���ߠ���
��7A� ��u?[���?�)>���DB�Lo1.]�<��l�����썲[�! �z�$��X�{c	�hFH������ʂ�����2����U��.��)��z���[7�D��6~�7pb΂L����
(m��띖�#J��>@����� φ�D>����%@��t�5�KF����|�2=�ܓ�O.,vT��N�L�����x#���q��q � ��<�rߖ��^#&���e$�̷tO(��3Qy��o�/��ơdh`�0$�R?�f�������\����M�jθ�l��:ޠw^���
���� ��E7��LDZ�&��v��jS1츜�#�m��.8���`���%�v�bտ�ECؽN���1ȸ�*�n|nP`�����c�%n����m��C�;8��}Ix!e��;.V��c$��� �T���*2m�DG�A����;'�=�1u�Y!��8$:.dEޝcxh��������~�]e{3�T�=�^��<a�y�tZxB����E�Zi�2������VOĔW�AD �K�8�$�|�ŕ����B�߮�_����2y<my�����oͫ.{I$x�B,�V�	{����>ZW��:�l��.�a͢}�%O���fy �e�χm?٦|����aᗴ���kAՕ�~��2TH'ʺCN��*r�Ǜ�;
%��T�6��C��f�+��ſ�����l3@�4y)7�m�{����tބY��M�L���av��:1�E໡tHn{�h k��`�K@�_�o*Ú��H�ܴ�\��XF���IBhqNe�^�n{?3��C�n/lڟ���E�ž7
��E�%kj�i|��S��� 
�؞��~%ԅ-$��Qa�\�Q�iO�fO��J�P�ȉX�bgg��i'����<�-����5�|�:Q}ɺ-�N����dko���Y�k�-�M��l�$`D��%�^L��B��Q�8 �4%����`��z�l��#���.�z�!q.䔕����V���t[����b~��D���ǘY�P#r�4lRbV�:f�a����tޖ7Ig�mI»�%5�@�P��?-ƪ1���ڊ!y����t�q�Ots����k"`[��D��*2��w�=�f=����{�X,]���8iS��tG�gfq�s
!$��$
-D��9�?ara��&J�}��a�|�0k��͡�{�F�'3�TI*7�U�u�<Bz+WI�+blI�|mgC�l*i�D��2v�uv\�3��E}���@��b�0��Ә� 5'�;��3����H	�(�C^��W8͢є��r�H�4��Ov�X�LY>��gAXM�)��v��s��*���&��2�~�ub��8��5�{ݲ�L��ԃ>&<t鍱�����S̥a�1qɞ�f����V�p�+6gs$)k :Ie�2ҔR�ꥍ_0�t2���.�����eZ�ȧ g״�"�(��I���N�����3�-*�R'��O��g0�iDx���`��AO�Nt5i.d�/4)Z{~�N�c_��e�XY�s�`U�b@s��9�z�%�ȥ7�I�h�%hu�:uw/r�M3}��U�k�C���̏L6h�U�slݜPX�OYa0�^����"��1�fp����Ľ�V`#JYC��<�ۘW���%XɄ��d��q;�-��Ix�vy.=f��
wb�*�p���I�]�/z�6���X�t}���ꗻTɑ}���z9d
j�a��o�ݽ3Fo�@:��h���-8��V)��$�W
U>��5�L��:��WW����\P��
_�3�'֎ɟ� v���@�Ǡ�8��\�]pVW1�9|�~�(|�0l�ebr�*8�% ��-��{�s���$8%\K�PB�%�1Z�$h�?��%��(�s� *�\�~[��8���`��F�OS���G:l�o�qKd�o�~�i`>_������<1�To���ߤ~�*UO�a�?�����z��T>��RyI�r�Q �"�x�l�3F����Ck{���r����
8aaU����&0���RMuc|G�������몳 _�e�k��������/X��T�Ǭ�����e{���	c}�C�1pWZ��O�Q�~spф�`�z����nݲ����Sq:>f�Z�5>�C"6}W�hן=�Sg\/��p��#����K��8ܻ	�pG9�<
'i�]��t������q�h>�)4<�!m��_�Y���I�}�Z&�W�gC�P	�+z#%⬸��8��õGh�3ç��f���M$��2[�*�c&%�M5Sk(�CX���i�tz��؛��O|�X�w��r��
𧤦z�������c���6;Tx��z����7�U��l'2P�ɠj��]�]�	�5�s�i�Y-?k)��Wxŵ]�K��eJ�4]Ph�%�+A�p�I�|.�x�PW�=���S�W2��A5���dׁ�!(�~zG&`�J��A2�����$>"�z�
f��\�؞�=��Y�9��\ޝ�
;jn�w_>"�ߘ(1cy}����<��0�sjq*�w߷�^�Bd�g�ZE'�MA
ӈ+�-v�����Q����ܿs�Mw�j4���II�æhN��YW�����̟�<�
X���z�0s`���T"���tt��I����ө�t�R����M\��H76Q����KG'�:�=2wv���?%o(h{~%���'����l���됖�X֥���ĉ�A
F[�� ;��a��Q�;��ƹ��������y��abh���o����#=N�K��AKU|Q��Z;T1�������f���>��4.����^��a�� ��z��}��r]�|����h�Ǣ�[����pLM�� N���7`����C$��t�\���GN�{u��(��7�`�X�:v�X'U;��]���'C��,O9��P��D1��80��ۣ3q'���$�J,������ˊ�kL�*�����;���as;	�0d:�ۉ<-��*iȍ�vBѓO��ʔs��L^�o�R����2��S��f�b�nP�������;I����5o1�1x�����Pn5��&�gl��,��32e�x{��zQڃ��S:̇�����? ���(�魉p9�����IS,�W��ג��⊏�	�a�Դ�e��͒�l��fP^��|I��^��L����+b�h�������q��CK����s��v'��=\�"�r�(�����K4�-sV8"�yD�mK�t�?6^��Ș �S���f��e�il����`���I+�!�
�����u�hU��w�?#�3���j�#{�1�XN�#���UKRzE��8!�"�0�n��w�K�=��CΪ��f<s�.��4#k\`i���&6[�e����e��v��}º68Qλ��ͬ�a�*v_i�����K�)�_V��~t�ISle  �pQ�#���Kd��g�Z�b=�0�R�N�d��1"���V|�EʼlP�Z��<�ٛ�ӲR����d��mC�D�^��-��K�!��|Z�V:l�)]�̧�sR�Xpb(�
�qZC���F"�jL��@0�X�@T�9�~�t.RK$�iϐ`G��H��n+QK�l��wȦn��J,4��	��N�g�."`�&{�iԳ>4���o&�up�뭗�C"XH��Rɒ�����m��������E�Zms��A�YIdQ�H/�|վ�|��f��"Պ7{Gֆ��Z��/u�Ī�բ��f�x�a����.����.�Վ���y����a0�.�^���[ӝ��o�5Mu����9?��[�ڰW9�^�q��vPig���h�Ϡ����*ҁ����ʦ���0P<=9=P|�Oۄ"�	�^���J! ��L�]	�1$��i��F\�"�gP�Nx)���Y���d1��Za�ZP(�)D [83�Sֽ}�%��쿰4��!����Ϛ��`%���8�6vz�t���(��~J���� �]r=6�M�'%X��-���@���cjH�o��� 4�j��fhA]�f,@���m�*�����=T��~�-u5'!�6Z/�jM�ˤ��u�px�����&S��Iڵ�}�8jy�7��A��h����p�`��:�Bksg�s�⏞)�Ihj�De��&B�e����)8$�*����\�<@�O���@׫la�g�'���"r�eڼ^�p��Y֣�'r�8�njKu�'��)A�9�)%���_*Tu�CU�9YFPQ��w�O �5�i����V��>�m�%�:���Wg�Ve��[���eiu���2���px�ð/���ي�n�N$Y%�5�۴o��ho����u�F_��N�oEߔ�+�{.+�]w"b�C�ށ��h=�G�9���y[E>�������7O&���eZ)AM)����}����	��s���V���۶����7h)��{4�G�<$�-�'@f���O
�Z�O�U��]��>f��Ǡ�1D䐚��i��%1N䧉�]b���B�W������G�G�Ϫ�t�t�`��\زe�B�o���C)�ʣ+Z�P�e��0oz���9WVB�Hݞ��Y5��9dV���/�~ә�9���<X,S��.�h�v��k7?tB�m�n��8�o����B������$^�	�靼wK��e�ͭb��OG�,R��`�NП*,����P.^-$L/���˱��G;D�5�;�P���:�~&�$q�`����[���@��w�̿|���K�,��8���rm���GB Ϗ_����Ѐ�̔�*��;nT�J6���ٌ5�w�VI�NhNt\�m@��!l�\f��%���y�����mA�0b��c!G�Jw�+,9X���a�n2S��u��&�(��!zW��"c��59�*�ſ�#C�� ���*pJ�U 0�%�|�no%Xi����������tI`�

�܅Әʮ�U�����S�n�K�t5T��9#�jv����qh�`����b}\�:�Y$��W�{<{�8
��DGj΃��_�#@a�2�W	�l��
�����Y��u�,��@��;O��c��I ѭY���;�/(�bVr ����2U��8p4P�_#��;: ����ɐ�\���Ԑ�r������uOSS���]*xĿz��*�C�G�{jb2���j��]^0��9a% 8�/'^{{��MUH2�E����R�e���i���?[��yp��|F1\N�0hq��R���U?�}o�e�t�P���S~8�K�?�J((A�F�cvt��h`����j$=F`%@X+�I�sgU��\cm�ApA7�Nވ�^!�y�*[x��~C���5:[1��uC^J��y6�?�-��@�	�/o!;���)��X�̪;���I}���)�̦'�+��,#)�+N&
�ur�d_0��ȹ��L�_����T���B�����;�ݯ���aj�.��Ghp�����!��@zr��>Jį|���QQ�7��:��88��oC󷇜t��O�����Q��6R�"�&��v�a���ԉ�اoWY�n�
�����ay�"a��}��rC��<���q�Bk�>ӏK��^����5Y���[6�c}|�>C��eV�ݩ�k
���B.t� �����s��a�T����ձ�^��ݞ��ڍzx�F�h�B��85���8,4��5탧�ŀ�Б������C�	�72�!)�j��j���՚Nd��m���voG�=YW�ecd9{26zv[��(�Ă!$������l�v��pW|~|�Zi��c���5\f��f*�������&7�;��^i�?�g��S?z��Ɯ��d �y���qݮ�i>a���pV/��e�#{���s�F����>fYNZUL����ԛ��\�
T�F�)Ș�10��U���\�beI��e[M�^\���i$5�,����,��q�.��;�䧔��Ә�'���K�.�v�dU�>��I���@Oq����߭Y�v�׮���'{9�(f<6��Ǯ�&�(ܒ�\�faE�ie�xN���
��K��e�:���n����>�V�v]��Qʅ���6v�⾹�r�wC-v, N-<S�E3W~��7�hщ�!��귆�����#�K��;g�B�UTy���:T�)+u�i���c^�nHeь��)�E{���dK�a��� �B.���So��SW���ӆ�����гHQ�iA{ĳD�j����6�ϴ*�zFN��f��>��1$�:���e�$�L�%��c;a�L�/���3n�(z�D	_P�аu���T6����0��M;RR�����xԭͬ��a�T�J�{�@t"Eڜo�t#byJL?�$�0|�����&�h��^�_�)�i´���m�Y!�O� FϾ%s��j	�4\��|8��jJ���CwY	寻��AX�(�y��=��$V�zR�Y_�7}�k�UA��ȲsW�<LTҟq���*�Od�S��U����@)�6�NY���CԻ�.�����?@�ZapzU�$�-��k٫6��!����:������)^<�eI��)��L\�J��$"4jfe�h�I4a�g�g��/�X��	���o�bs8�yP�n�^�ړ��]V���q�_�����C�׮COM��th O^�Z��&yn��U�,�b�ʯr.��`��:~�����Y>�޷?:KWt�]Cm�V}Up�
AC$h�t��[dk���*r"���PW+�"�L��T�<LOPe�<�Ө� �Si��8ko�Z���8�T���;�pn��J���s�G)���VHܮ��3��2$������Wa��Q�����M���](m���0=�ViÄ I�#�l�,�f����o��i�P�򥓮�@�T�!Y	Y�E2�[ڈێ�)T3|��C��*!8f�]"P��Ò��?�Lz&f&'ִK�r��c��f����|"��cSlv_fA�1XG?������h�Sm�ÿ��N�A�c�˳��<4�[�-6��㠏1}6�x8���j��p�}�ٽ.����a��B,S,�nc��j���r(9�5mg$��-)"Z�p�^q����*��`> I�\���+$�fD{&�|�WZ~zɳ�j�H��F���`a<��c~G�h��}jF�Ea�#Fz���4���e��BXAd=<{�7 3(�E��뾀���F���z��$!��9�=���D�����t�K��%�;��GP�	��L��3�ܝ�~ 3`��8����xM�tC?R��,楑���F�%f��ҍ��BI+�\������b�i�t�D)�V��bm6� {�a��յ�$a�
��6M�'��+�-wٗfp�#�Pu�v��G�\���n� �.ܱ�e6��-���u��A�Hk�е��w~
ă>�G@�����t��m�-S��U�k��ա�;GWv��)��=Xnˁ�rWh����ZcL*��7Ł��	�o/�N��N��5Vha���7*ն>�N�H�ކ-�����U��N0B����Q �
~&��d��k�*zr��Ѕ�v��|�>�l0X�s��!Z���=G1ff��䖚ᑗE����[B��J�b��:���æD�<*L^n����/u�w�����]���@j#�BOңLW�dI�4\����j��Sz�	��/$Ho�$�ω���d�^Ie��� }�u�wM�e�K�ue��~�h{��oލv�4�ZR��t6��gjBǻ����,�=A���������Ԓ�B�ȇ�ʌT-���t�aweiÆly�
G��)�Ol�i�@�� ������T��4X�E#���QI�ǥ�!|V��ڟʢP��6��դ+}�W�"j��m��6Y�܆$#G|��(BTG�TN*n#�ݜo�~h��F�T~�����{Y}U%��Troq�N� ��>�A�G�$R�,Q6`�@�w�C�y��$;� *��q���}�uVۆ�݇����eIЬ�!1/��V8Ƚ�N4�NŦ�;�^/BO�V��J���B��#L�*B��|��8172��&�ic��/��~KCHn晵�B	��p��)��6��x�X�}�bu��׫�_AD��� �EcwRe%,�g�糤ƨ�w-�I})}��HB�t������;ܝ�s��N�Na����1hƆPx��}��+0��`E}��=��W�Jt����M��X�Cq�9=��y*B�@u�o���{	��/_U�E���>�ɝ���^}5�w�!/�3B'(�eC���)w�zG����$���A�I�-Ѿ�9�"E�I��eo���q����2�Fԡ�ל��3��ʝu�s��(�)�R�v�WSq��־2�ҲY��O\y�_>ӪT�2R�l$���R6�������^�HJ*���L�)�8s�O�q��a��5����c�|�E���(��cŸ��ZV.vDn��j7?T#tQ�Hi�~�'�H_�}��
J�?m��rܭ���`Q(��eB��^�+@�5�h�&<�k�}&6�gm�g|rNYY���u�g%�V�7�A�Ԭ�|�ڏ��URn�z�%��y�S�j�*�J`,�mO-f.��+���x4…Qץ�}W��*��iwD_��ރ���i\r�Ժ����׳@��c4Z���
)Y��+_b��#r+`����a掯=/|��G9Yv�kmT��Z�ֱ�JX�p ���$'��r���2�Fi�i�vlIxFm#9�_O�����k�q�6��evJo���eu��50[<*c.��B�H�)I8���j�Ն�N��`7n�de�3�?s�n�o8$6�������?��H�h��s&�Rrl߫� aIڳ�O�����_�QH[������jU��v�F���T�R�:x*O{�Գ�����t���X�Q�6��ե澓����t��}�a*�����J��`G9�)�;|���!* �tU܋�E��΅���_�C-s*����3�g������7	̓ЎǨh�ρ�R�/p�U;�(�#��v���;A�Gb���=���Q�i�{�Q�$Z��&���3��{h�3܏�d�jq�'�0)�<�[��΁��2E^Qc���Y���;��F�$���IqD��~��09�+t���^R쟾��B7Q�P�f�xH�t�%eў:��T_i��"Ux���	C�;�ꯕ��/�i���?���h����K�!ex�䰆�O}��g�m�޴�5���2d�^�A��=�s]��hF��4�I