��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&��n?��1ů��> K�-� �&�T�Ek/ֆ�\�놭5�DꢘP���+L+X�4��J��#�0�8���������l��jT��+�(���������6�MC!D�;�m�퓊D@v_p��䙋ⲝ��C_�6�Ռ��#�� ���	RD�4D��畓7���vn�H���0���fX����4 �CS�C`{��;�L����li��� y+����FD�p"��]���y��R��K�({� .؜M�������	^5���ɋ��&���&�@*���
e�� �t+���
_6��O<��7f�M��u���m(MrN����z�jL���@T`��M3��c�uQ�Y���%�dD���,�~^���y@Ga��(����C����	��G�86�S$��ɳT�ز8���:r��/y�[ݦڍ#A�����i�&<nU��<[5)�Z�-Ĭv���0t���d���"_���:�'-��d��*��q����_d�y�N-��~";#��������Y��؆���	6ZJnԷW��έ$Y�K�?�4���L�w�Wmiɶ��Y�?jx#*�i���F�m�E����O6T>]i�_�9;�!(��kH7�OS��_��[-M�((��lO�s�$�g�x7`��ZV�E���F��,9�j	@���]}<�ahb5~ãdl&I^�	v����-�@�@���	��!��d��`j[Q��� r��;f�i�.�m+UH7��/OV��c��������l��i��M��*'��?���G� SK�M��H?�7�|��}qz)(Mx�(��ўӈ,X�߸���n#la��E̺�cRe	�cz��-�p��N_�:tB��/��>�[2�Sn���ۓ`:�iLX�>ZM��<
�Vu\N/d_���ۧi�Û϶����a]�������A`Wؖ��>Hu�W}$/])b3ؾ�ܙ�9���}�!n�!�
�^6����9�Co�(���0�X�%�<z��H�����&ꗄ�5�w5��}��oL�J�ϭ����M<���i�ؠ~#�Z�R��U�>�6�՞ŷ5dȿl�Jj�~v����EA��[�bsҁ��/�K]�4��<:(�*�'�OC���/�/St�e:qyeꚃ�T�&�\biM�վt�,�
qdj�8L7�qt�J!�&w׌�6���R�3�����0�H��1r�n�)�I|8ȩP$:��i.`F��2�������rw���W
���L�X2	�n�K|!�<_e�1�)�L��.L��*�D���l`Γ)`��3,q�T�kc��2��u�J>X��]���Tǝ�c�5i�*��b'O"L�5@	�� 9;����)Z_N�z`���}�9����m�D|m��
EЏ�9���!fF�a������,�Y˨����>�VmP;Yjp�A=z8�m��Pp8����Y��Xd_��P��M��2qvx�y(�n���p',��*$R4�BH`����=�Z{�
��(�v�I�:=�Y��])�iREf<�+F��0[�rZ|Va^!Tы�������tڋ^�T|�)�G-��m�b��;9Q�Bu�ި����^�,ji�F��of�01��"n��6t3�q����%Kٟ|��o��N��M�J���Y�E�74�^�<	S�mIr�f���C���Z�Ŭ�ͷ�h;�ӼW��r���F��s�a$;��GNq9�����ߏ?���:�[�&�����?2��e�!v�
��6��_�"Sv����s�����dd��T��6�1Z5���:Io:��D(��c`{�|��#muAL��4At�/�߭�;9E�e]y�qlF7�DJu'xi���������e��D��|P#l�����<�	���ž?G��Fd����Mj�'w5[�@J��j�?����:`�\�t��[;�z����CG1v�Ƿ����4�/�Z�-:Q�1�D�j�S�	T����Vj� ~�Ҁp)�0�z�A%�.��̫��:�|+���ԧt�W���;v����i=�z����)����������=�/�+�O"��rM۫\����Ґ~{C�՗�e��ML?;�~x�`�Ra��3�lWP6��z�8�
\��ٚ��j����R��2�I���ʕy��r�X�%Dv>cǃ&�)��]�q��o.�]�������&���}�ܱ ��1�y_օ�Zf���g��P0���yC@���I"  ���S�:��d����C?�R���ӽ�kz��&��LA��r+M�%'N���D �[O9i��5Z�t�^]��l�o~��U�����|W�FF�4��8�<�	�����
8[Rh^WčXg}�������q��kay��4��]).F8�h�A����x���jZ��Z+Fa'��m�]j%�ĭ�ƾڃ0��O�]�ʶ���-���Q
����}+��j>f����G�� ��]�4gܓ����o਺��mV����5�&×��N���Ý�{9C[��DV�3j��֨;�7��s�2��l�eƁK��7�����	�g�	�$���������5�V/�zTZ�s��Ȫ,Zdl��H�>��[o-�Y����,4��iڪ��7�8cncg�{ρֱ����X���d �6q�rl��_Y[2��1V��c�JZ���榃��=�5:�P�鶤H�^AB��@ww��Y9���l`�N�����R�3DK�Z#��k�-q��a�);3��r;��Y��,9���h��Y�u��$`5����dZ�jPŝ���)I���\4�Ԋ+r��+bvQ]&����kIN��S#�A>�
s�SM��3o��{�cm�Jw�I�LM5�WK����[ ��NH��;�\M�@���X���A��.Ֆ��-P#d�Q��'d=�t��u�^�c&7�ā�7|�G�]���u�����ք;�n��KJ�nbc�"&�i1��u�բ�=�;#L�wX�� �L�8J�;>�A���q9\6j��!Z��yx�1���"KGk<����s���L�,�r�1�h2횮и�� #�&Zum+L�����c��sܕ����Y.�tݒ6�������5�uZY/�ϡĎ��,�U_h�L��@��R4s]9�@a��%��ɳu}J���i_�����B��w58:�Θ��r����LT�_��Y����^c������]��%�0�7�s7!N��%:0��g�.�m��������h ��7����Hq{�������յl�(�ݨ7���0;����~��d�HZ�j�W�����K0�8���<�Y���]��]�����s���`�<���wJ3��f|���{�{&#j�:מ2��|L��ު�/����MI�[Q�}���`_�P; �����*�*#�Z�;_@Ih�B{��>����5;�Eƅ�Zo���������s����R��ӯ�������� ��B��YT�X�⦣~