��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&��n?��1ů��> K�-� �&�T�Ek/ֆ�\�놭5�DꢘP���+L+X�4��J��#�0�8���������l��jT��+�(���������6�MC!D�;�m�퓊D@v_p��䙋ⲝ��C_�6�Ռ��#�� ���	RD�4D��畓7���vn�H���0���fX����4 �CS�C`{��;�L����li��� y+����FD�p"��]���y��R��K�({� .؜M�������	^5���ɋ��&���&�@*���
e�� �t+���
_6��O<��7f�M��u���m(MrN����z�jL���@T`��M3��c�uQ�Y���%�dD���,�~^���y@Ga��(����C����	��G�86�S$��ɳT�ز8���:r��/y�[ݦڍ#A�����i�&<nU��<[5)�Z�-Ĭv���0t���d���"_���:�'-��d��*��q����_d�y�N-��~";#��������Y��؆���	6ZJnԷW��έ$Y�K�?�4���L�w�Wmiɶ��Y�?jx#*�i���F�m�E����O6T>]i�_�9;�!(��kH7�OS��_��[-M�((��lO�s�$�g�x7`��ZV�E���F��,9�j	@���]}<�ahb5~ãdl&I^�	v����-�@�@���	��!��d��`j[Q��� r��;f�i�.�m+UH7��/OV��c��������l��i��M��*'��?���G� SKٜ¬'�Wx�R�4{�ŲFRe����v2�	��t; i�k	�7
U�<���<�l�r�pV��$b����}/L��&�q��!�}��r�i�+׮+(s@�����K]>*D��E5�R�b�g�������y1��	ET��r'7�*��l<$�!�O��n���^��rnLzŉa�c9�=�m2�3�QG@/f�mwV�5v%k�g�1�m�H1�D��(�ɼ��n���4��s�6�����O)�"3��OZ�,��.�p�F�qׁN$"x����F��I�Po��������Qe�S��������?j��7�ˋQʽE�Ե�h�)���kb�PEO�����$���u��(Ze}$�&y
�O����D�-��Y��!POOB�.}BW�K��Ü���`�f��
��L���fD�
T���*ܜ����.���|>�eu�5���=��J0;�=�h^Wp�qiĦ6p�gXDA�i�,��۝��j=T*D��(�O���sI���Q�U/E'�t��z�0ѝE8[�^@��ҦP8�L��)��$���/cC�����q�� �$'C�<��.3��s:�B������T�����8�*���<���Q%���E�vJ�>�B����X���:���n!�>�h�|5�T��t����g�!����E�`�i���1Y]��fY]?�7�_,:#�\?]XP�ߺ�!�O��ַ<�m� {A��N:�57_�^7�uX�+P����}��w|�bdE�E�N3E�G�����S�h���缃����������~&��vڷj'��K�ɟ^�$�yS�	���1�%0��:��B����9�|6-o63{����lk@�����u��}V$ڰ���ݞ�.��o"1I�v�K�Ws�3��a��.1�	�ݰ������2;q�֝˹��ؚB�'jJ*�S��D�FzrPO���C��>��H�L�-Kv3��pQ��Ps���N=�B��Ti�,�z$Zi3DL�iԜ"c�U�$:��8�T�7�zb�nx�h9��ی��͔��~"������(�.i͹?��lY�֡�G����Q��$��G�Z�ӘFT� /�R[���1K��U�4���&����Ogk������ԏr\���G���������r��� ��R�����R��>be����+����Z0���V)�f�����"���5�DJ��H��0��1�{��܊>|$*Y�b��?����,�a?D1##�Z^o�Yp��g恘p���Yj�F��_�:�P�y;�"����ҼXg��ㆊk�OF��"�e��<m
|�_�x)c�y�6s�O������W��zPə�*=��J���`5�M����ϫ�^9�Ε�ͬN���#���M�k������x�[�$�����}C)xi! ���6Sk�<�I�g���MĲ>#����ˎ�'�o�?;�\̧HR� 4g(�om_���L�k7iE|�f��!��WI�n�?�cfJ��f|rH���c��<�A�1���i����4��܌�Λ\2�MDK��='��Uú�>BR���0@)�CG��
�	�`B�$`��Kqe����$7)��o
e1҉�f��tqk:������\<��.yuu9�v[�4l���C��F�Ǯ���n���I���\4��٬���6�9� �?�xO�)=
��B��l~����i���?�g��Ei���=�¸g�_��Z���?�����u�ˬ����鷔nw�)���vK�0�0�X�Ic<_�M�o�x`�V����6k+�7�����j����+V��C�;}�X8|d����
#V~v���m/t��+���X��h�D��ʙ�ȌիQp�5Y��P��#sy����vɚ��{��͖�J���2'�eg���4�HR��\���S����{�;���:j��8�D6I�(ITj�O���żF��w8bּ
�ќ(@��`����'�c�Z��1��}�
���֭��h�37�$�cW�<��.+��7��QL �o�̐b�D3[��
M��:��1_a]TF�#Cy�zv�PM�#�'>���[��I��;?Ү���5ZdB E?�K��тI�WI���;�CO��|j��cՁ��f��eӧ��ZՑ��$D�lϜ7G>����ch7�s��q/$�6c�d`�$	�8�+x���Ko���t��=�ߑc�qŶ☃�;�s�"Z�Q.���'���ՠC�R��b/A�j| {�k�n�׋չ��ق>�F�$!w?'����p6/�tWg�Ɍ|��@�Iq��f�g��/�PP�/X.,lH'6z��FK�iO�B����Ó�!���dx��,xv��mBI�U�Y^��b����MP�ʳ������Y�8᎜���W���]Z�,�k���;O5���{ʓ�M� �Ztn�3�5���+�T�w�Y�*������(����R}"���4�%�4�bm!5*���Z��N��L��b�� pA%꼤G���K{�^ah�j8D{^�箇�}+N�ГkhW��윯���`'���YŐp�݆���>�k��n����\>U�`ܧ��������V���i�(xO�BE.D�WD������˘��sf�o>��+�z�hC��1o���=E�Ԙ���9!Ք|�x�E~�Go{�1��s�X���9������+?zm���<�Rܚ�>%Q;�+/��϶��k-W�Ӯ��=�%�a�����]��h n#�}��7�#��4��JO�=q0�;F��5���=��U�I��**�O)�y�in��^���,����k����@$c˒��I�_1ȍxyw.�ޫ�)��^��FW�$
9���k�*��Uܘجq���`�"&�.o�]����{�<�2��^V�g�l���8��:�a(�3?��4[0�݈^�R�� `�����_��-{�'t�懆�v��;Z9��I7����0���D� G��@Ƕ��mu���JV��]�K�{kq�?�f�{-��H�ɱ6�`�G(�Y�=R3ŵ�s+��v��j�K��� dr����e���{��䙎`� ,|���[W�װ�Qn�Ӧ Mhr:�y�\z?�3P ���%0��f-�wgƌ�@^���;���C\J�>��A,ڀi���H.Plg$>�S����kMԅZɷ�Y��>�Oˁ�-�˽�v�P<d���py��}�+������n�E(�����8"�hV��w�|�Ѯ�"G�B�O���<Գ`L����`o:���x�jG�\�X�:�* ��Jn���~�o8�$K^O��C�).h2@I���1Ep�s;�8J�'s-ox���9�v;��A\��
�/ˌ���6��ά������Aq=nP�?Ǽ��\��vˑ��F����$Q���e�-�#����<�p�Ӫn$���G��e]�H����zHH� ����|:8
]Wyy��j�S�@3* �$�b��� ������*�g�L]1Yx���~��
/�r]7�6p�*N���s�������vU�Kl�,��K{!���®8�3<�@���x󨴳!#���ŝLBن�A�M
~��
D$����Ŝ�A��T�=�go��ey�������(��;v?�K��Ǧ�=':�b��h�ϻ�4�������+�n!
�e�W����+�E�S��/f��~��$4��!NL*�a�1�0�Z���,�"*B�{��x���R��%B��_�p8�6F���3�w�M
a4���Y�Ǳ����&� e�M�B]��Ñ�c����roM�����, _��
�=V�r�yv��ҡ�(Gl���7�V������p�hV�-�}e��a{�̬δܠ_)��q,&���Y��#��m��g�wA�<�k�0+�7(������Fo���PO��Ŗ]��R����+�X��GG����` K��Ȟ�a�k!X��(���cPt�ChNQţ:@V�g�J�7���c¤"�-�����HX�'�h�q%O+��U˸�7b�F`�����Y���eT0�y�r��V�T�D��i���$��K�Y߹Dj;%;��&%U �,p��m��
��F�Um�������q7��AQ~bڤ��ka
��!�Ğ���
��"K�������l��>^���?�?��0�U�*�WM�L$�!���<��EW8h쨵T���4�6$���@�+mA����������{}#��K3Ոt.�Wmih��b�+�A�С��%��A=�A_�Q�[��B�b���mK_I��$��Z�"�!�"h���v�`t���Ny #��"��(@�hM���2s.`�����}�t9B!� o�U;���Kw�"��u�A���R����{�ݿ��Ȅ*�M`�7\��M,�ẞC���J��\�ڞ&�]&T�L�`Ӭ���Aj�x^#䭼�ϴ��=c�Ƃ�ܵ���1�Z������:�R&,�B�A����S���N	gƥ;Y�Yf�>�Fl��	�z�a���E��K�?;�l��o�N���L)iD	�t\���w�ԙp "B��rA��J��>t���0�[&���*g�^�����䓐uT���.C|��?��Nޞ�sC��OR��,kc��O�\̀Ƥ2	}�:{��H�A`���;'�87�sǴ�e���4�b3̥��Ǝ���Y���Y���'�� M�v�_ ����5�;$�@�u��d�8���G������|` 1�_i.;֝��}�b�a�xE���w��Z���������ص濭bF�� �Wޔd �G�N!�X�Z�wK4� J0��m�պz��K*j�܆V�5��d�aM��d�,�*����?A?��7^����)�;���"��f�;h�	�
.^~��/Z���0�:�/��>�B�Yӑz����7~Y��=�Q�J\��Ώ�%���yw�\�:Q�	Z�]Rɵύ�q�q h�}�״��N�U��I;X�<��Iy���{�~ǎ�?�^���>k	K'�X�s��:�Y��l��m��^���	�
�W<3y��ӴMp�]�>[��GY���ߨ�xC�>��(���l�e�t�|ąo����؃�hn
f���=i΂_r�P�y��y��VGl	���C!3ԑ�������.:�wq���Cǹ��w�pH�;w�ix���=N�ҏs�82��#�zQ�\�&�|,�'�k_�T
�3��,�0��F�Po�S