��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&��n?��1ů��> K�-� �&�T�Ek/ֆ�\�놭5�DꢘP���+L+X�4��J��#�0�8���������l��jT��+�(���������6�MC!D�;�m�퓊D@v_p��䙋ⲝ��C_�6�Ռ��#�� ���	RD�4D��畓7���vn�H���0���fX����4 �CS�C`{��;�L����li��� y+����FD�p"��]���y��R��K�({� .؜M�������	^5���ɋ��&���&�@*���
e�� �t+���
_6��O<��7f�M��u���m(MrN����z�jL���@T`��M3��c�uQ�Y���%�dD���,�~^���y@Ga��(����C����	��G�86�S$��ɳT�ز8���:r��/y�[ݦڍ#A�����i�&<nU��<[5)�Z�-Ĭv���0t���d���"_���:�'-��d��*��q����_d�y�N-��~";#��������Y��؆���	6ZJnԷW��έ$Y�K�?�4���L�w�Wmiɶ��Y�?jx#*�i���F�m�E����O6T>]i�_�9;�!(��kH7�OS��_��[-M�((��lO�s�$�g�x7`��ZV�E���F��,9�j	@���]}<�ahb5~ãdl&I^�	v����-�@�@���	��!��d��`j[Q��� r��;f�i�.�m+UH7��/OV��c��������l��i��M��*'��?���G� SK�M��H?�מqT'J,!A�h���'� D��G�T�>��tw�ܻ��l.pRu\7�V-�T�V���CS@�ewf���H�*�cwl�H��ϋ��#�`IY�k����_��U�A#���z\�yz�~�cٽ�bl����S�&+s#�V��%��ӧ'A�N��qT�7a�t��$d��]sH8�G�?����i��i6�ˋKl<�O/���	w�C��:�D��]�l9�ތ�G6���Ccyg9m��<%���o�m:|0�\)!�)�2�*�y�e�M��%����� w�Y�.���,���E�ٗ��N�*��O�zP�i8:³��v�\ݏ*�P�?���`�l��F-U=7�g���w��ȩ��$���"5��!������{Kh��������k�$V,[No�"a�K��H��c&W���Xu3ѳ����i�uI(of���p4<t�Xzf��4p-h��,����<��W%P�)�������c�%w]������"� �ۭ��9�[�Z_���K���N��� �{����Z�@���k}]�s�yR��݋}�k���/���7�&�<�V�0��dG�z}af��5#8��N1�M ��Tl}JĖ�B�	�}E�}�A�	K����D'�R�g��=	������+a������%s,^m�����Ԝ>�m�����?��/ ��#]>؊uN�\���0}�ڇ�T���cj~9�I/g�~0��1���'`p�4��w�:�)�W�M�^�p�r8�^�XO�>j�̫h��BZ�T:�x��z���Ρg��ldQ��q�!\�_p�,�>���T!��P$cx׾8�(�ct��Ζ�6���yV[�WQ�;E�p4إ�d�jϊ�"$F3����]���X$�к��#p�Ԧ�ǘ�����j�s��Ղ[%N�~:�Ls��-����Q����c��Nx�qW�k���x��4��:6��|��H�������ۦ���'q����Y�5q����/����AŜ�y���=$ g%��'��Io�%�gj�fS�rF�q�O���)��z���Xff�⟩KG�/�}	Z�4��|ׄITˢq{}M9�K�Bx~s* ���~%�m5������7w�Ɇ�����+xD�ͥ�)/G-�+��{���e�7����"I��U��MIIT�/T���`���|�ƞ�o����wܪ8XRp�U��3���ҳJ$����A���Ro� ҬU��u;��f.s'cY-��%����P�2�#��x�\��0�oae���YO��!�6�9����g|#�O�m��M�=9�NT0�Ɏ��]�P68uT��M�)���@<|��+��Y,_���Ж�Z��_��@����J�qL{�} ���/Ʉ'��6?�P��V���a�\��#�K)�I �r�!����٩F�����SS�_���"&�zRf�xL��y ݗ����v>�0>��h�R� L��e�����I�9����!����\M�L��p\�p`z����@6u<ź��j{��7&���<�.C��v>ʰ�����B�b��#�Of��l�1�q�fu}E�x���Oۉ����ʧ�{�^�ю.��l��X�E���H͎G-�[��!��4[�;���1������n/X��B��U���Y`51��P,�m5�ۖ���.�H*�G/s�W-"SnezPhǽ�,��c� ����o���
H)�(j�V!�������>0��?EF��E����-��Tʤ���|�U>��$�G��_����$�w����d��&�({�38D�����4���٩ܻ���L_�V��G����N���sIټE7��ϙ[�ktY��.�S"k� ���\y�������*���T�Ƚ���G�CK�!�څx����v���3�?Ѹ�7�M�q'�ـ�~DZ�FyP�u�9���k�޴21!�f��ZN�q0�=j��",�����k�|0X}����m ٣$�R"|��gZ��Ȁ��ٱ����¹����}�Jl����ЈD�b
"�4S�q�Cו�B����?��b놾���I�E� ģaMY��Ġ)jc���3Ԋ�<�p�'"�s5U��F��woUR5�#�U@��a��o��\�-pzH��9�Y����3��;Ј��h��f�8E�Ī|nlggFp���d���謯c�S9� (X��G|��s^@���<�l�c��YrW����I�45��4�m��n	��fG;���:�.凨�Y 2�]�a)my�o�-�b��:�iF���X,��M���^f[�W��g�RN42&�M�z��8)5"Ն��n\�X0�9��{^YGG��8dڇ�}	�F��/��Si�GJS��^N���׭oBN�5F�Z��t�$W�j�K��%�1��� p'�vٿ?H�Uw�]����JF�_,��_�ާy'�1J���]`���^���F�HYq7$��#Q= �a�>q�V��{���Kɭ��YZRO���&W�OEed!SH�jn��Mh��"���D���ɜ�P�F�
b�ca^�x��=!G�= �0z՟*ի���6�)N���9�U��,Gw��%㽛����u�%�j�8|4�l�����^(��q���h�ӯ�c����F�#�\��Ν�T[\/�����X����L��z�o�d�P�3�h�()��͐M�8U	�~�=�ǡBWR��.�K{:jb3��29��Q*~R�'G�����q����G[P���R05���mI��{U�s�d�j�7M�z��D� e���!����ʉ�j����_g.�Wna��ĉ�3�����V�����Ԃ}�l�?�c'xI�wa�՞��k�.ި���y���H�[&�M�&��ɰiöɓX����¶?�Q���)�zg����*4���4V[�ِ��O9�b�O?:/�I$��Y�����b��3�۟۬8���K� 5���D斾�%,!�hĎ���h���ڭ.
�R�P�Y���o�@�v�D�a�}��U�"�c?(��3�H��m�tڒ�`�
�M�)J����}�^-�wk�찎��?�c�Q+����޹8��ʑ��>�;L���L1�ͼz�VI����g�"�C����?�<X]�������hy9�j�&*by)<F���Zq�r#�z\*6U�.���vr�����y�����W;,T���N� ��c<Q�eb4GK�m��$��ɑʣ��{yO��k�Q��B��k�-0�"��o�$��nD��ٿ��Gpr|nz���|Kd�)�<�v���7zӍJ�&��� 锟��C\Gn�O�������J�\,�UBqɰ�W)Ж�dل���(\A�XWP}��\Y��п! ��=m��GMn�FP�9��8�\Ʀ�f�y���{�Ϭ0 �/l�s_Th���)xzV�-��H�А`%�Ϟ�)Ù���2Ԝ-�l�'Q�v�~7��a�
�;��^(��}5�?�Z<$+�)�BUՖaX�\��n�c�D�̧�K�[8�8?p@�7���zz�ov����B��� Cg��u������@C_���yd'5�7\,�Iܻh柮<ގ�F~��8FI��8��jY>0
Ք�����V)ET�l,{������!oQ�4��J%��i;�m,���*'�%9l*�+|mF0�>�y�xJ�uN�Kц|�l��m~�8�v0{��b'��4����Sg}I2��]/�+�v(���eMw�s_�_�m�#�Iw��Ld��J��-�K&A6إD�.�u��wQ0�H֘ŘB�j�*I����8u `N�n��L��O*��%�-��)}�[c�n���;$w4�vd�K���Xm�ɫD��*�C�ܼ���+Z{w3PZSð��dNX􊳵P��,v�h2�S�c"�z�F>)��?��zAܔ�~�Q0�zDŖ����7e�+<�X�Y^igZ�u��YT	�����SߩQ�	��!kM�wwD¼|������i11�sC@#���.|"�U-���%D�O_��ݬ���tiAP�&)<��Ԉ�R��L�4���)#�;Z���<�|�`�7��ղ��b�N�.b�V���c�]e�,Hy��<�O�V�q�lpܙ�d�*W �7a�u=sޝ>�צ�C�c��>�A2@��v���^��(,9A�.�	.I��b�ܨ"O��ê���Wf���[}����:;���S���yw��%`%�}��o\�T�i�#x����Q�.�X�?�m�W�w�J�±�XbUyI#�v]���#�,^Z΀������s=�Z�β�d�n�p��|UH)�"��hO)�`��J��$a���E�ܧ��B4�I��kT5��n�#����`�.PC��+�q	�=8��b;�lV����&#mwʻ���w�?�P*�{Ȑ$s��u������W������Ѯ�c=�D��H<gm@.<�������� �v�|�"R�T���jӣ'w6�)�?�MZK��6)kIk�!e����7 ��31�l"��Z��t��+�l��'�qı����<���! .l�{]<z�=��OJ�fx�y{�����Bu�	C�D��� h��PC��ץ
 Tʧ��D�A7�
s�2r��K����zGv('�T)j�w.�����������U���&�G�3��Tvo+�A�Q��i����G�+F��;���:�l��r[����#�&�`������R�J���GQ��!��95�$�/����g�T(�����6���W�W��K)�Iԗ�"p&�㛛 joJ�k=֤Yq-��s��������F[�"?gf��I�d|��d=���T�K���[�2(�^I�+�m?P��"���af�W��[�O؆"��]�Q�]!��̪��+�HO���3�'�9�r��?P%�k��a]�4��i����A�ə�%n�z*��A��S���z��+� Q�A�94���s�W�H�����)~����_lw䦝di`��fq��T�����9ه�B�ߌ�F7U�۟�%�:"bNj��By��6��b�O��D�x�)9͔��.�kbA�_����<^��A��1�k���@�7D�w�b��)b�`�ֱ)��IE��4:��*%��g�81���>��T��lGNսw2�'�2�[>;u��`M�&�EW������1�-����EvQ�)�����7L؟M��6��Ӳ )�O�������t�����r�k��d�������ʟf%���6���{�}zx���|��\�?F�ʈ�:9�|�/����׾�̂����0"1�@���W�d;<���OBN�b�nd¿�5���}�z�D��0�u���o����S�_"�6���#g{���5����R�E.C�Ƒ����z���1�<T�[�R)���X<X��q.��m�$�s���NX�d�Tj�El(gg����ak :�M�����mmZǶ������j8��!2��
�*�B'�JtK 0�E��%���	쪻�A(��<��6��&����x�sYf�J��ˏ�j��`�6:��BE�J����7���s���қ����0�I����,��,X�l�-�&�&Eog����׽�ۺ����ݣ�]B9[g��M�k��MM��%��P9�Z�\���
v�v��Gpk��̬7�{N���Ǫ2��ğ�+���V�����wWK%S�$k�¤F�?��~��e����f�|�K�k��t�a�KĴU���#�ɲ��`��aX�]��M��EoSoR�L���㶱x`8۠7��|z�\�"�{s����IB�����*<��H(����C,�v�!��9�t~J�zP���o�SA��Yj��ɐ�.78�ϛ�T�1�7`�>q�Y�P�UA�U�+QZF�M���'|�+<��4'�&x[BH=D*��m_W����2�C񜫵��	�1������T\�(ɒp�i�C�O����&��[v���O�h>�n���.�U^����0�f��3�-���܊G�՛�9'����#���Qؘ� ��j�S�q �)	��W��xS�M�la�Ĵ�z
ݸ)�lnn�A�<Gп� �f�G���% ��BoJ��zPȕ$� !{7��������\xɥ"��*&�>~B��5��5*�ӵX�gd�B�Q��;���G�W���y�I��dT��,Z����D�ܮMg\sr�ɟ6H��55A
rD�Q��Pp��^��Q"P@�\�J8$/zN�F�v_̝t���!@��6���4���S2�p#ށ�N֊x.��Ĵ���~�0�0	�rv*p��������$�;5�2�X3�sB�1�R� ����i�����L�+�1}(���'���w~��p2o��e�6i�-E�b*6����&kW�L��kP�O�d�� Cᙵ����]퇭/ē�}�BZ6T,w׷��MI<�n���;�J|9}:�_��ݞM-�G�*�ty�����7:�E�G� о�d��A[]y�'IM�z�û�])�ě]C��3Y��Y��tx��&|�5�m�F&�!*X9 #�"K5(T���",��۷A?��F�J��JWn�/��8�
ύ���o&a2iL�"%�����@�{Z\:��t�����3h�hg�#�}�.�M��Z��sFs1�K� ����*Iw�����W�zՇ͉eJ¸���,8w����¦�;\a �ua�l�e�IZ�~����ť��ʯ�����E)���)���F냝J%e��x�M@)6]l�@�����;O�P?4И��S��*������n\!�K��"P����q�����x1<� M!�(i6^W��')��U�"D��:N���k}���H��`F�5�5Ĩ�1�'��-%;����%]��{��N�k:5�p�f61K\MĨ��>������1_��F�f�%�N�_�N��\^J������3GoC�tyҴ�$���Csm� �u]K��_�N�s{	��7W�o��f(�cS��J4&��sZ|b	*|דǙ�7[VhIw7^��Yz~��:���;"3m�- yJ�������ڪ].�u��Q�ᄦi(�ݢ�zZ^%u-��6�>�<[t�$�]ƱF��6x�� �Kܜ�
�^���%��"�R�\G�*��tz_�~�t�<�u�mJ-��dy��v���d�S��?�����J���)"Չ�7dw����Tuv3d�ӡŅȶ�:���/�g�������~lJ�L�IGℰ��KwEV1�gsF�p$���ni�*HX�M��n�\�M��Қ߳T�%G+ )���{��~�DoS��[��������\�&�	(������.�Z0����J�5S6�$�[Ym���FS
12�` ��d��Sg�~�X4̂@�*��]+(���?�<	>9�6��t�!��!o�5ڪt�#Ň�Y���0lY{�߫Q �֜���O�o�5_U��>8Ŋ��v)pW�� �E���?\Dc0�O=~��Q���u���ޮ���NvU�`���^�q�.��r��$! e+�H���Lŕ�!94��qx�"�	�\]��M�NJ[�|2�U�ڜn�����Hj�!�+����O22������E[FVA2��R�1���+�_�z�S��1vՔؠ�M����{�vx��[�K �_@��ٕ"��e�С���*s8\��+�ɼhPx҃R�'��G96B�Qd��*q��,��@1�����/�c�P[2�Q8^���3�O	��#+�uw}'��]u�@ϔ��$��Dz:����^�ج�[%�m�TA�3�,���ݹ���+���N�c4&sj)�?hefd�Ÿ'�֯�>��x�LvK���`����O{����'�ӓ����3b��[Va&���Etp>�O��#�i�I�����|�r�X�s�Fp(��j�8�"����#Sk`�j�<}}]d�`~���"A�rd	H���t�[O>6*۪��8E�M���oy�}��M@ZL;G1L?���MvMYKE��Ip�"J�Q_�I�;e�b��+pI@�ܧu��/8�3EӮ�i+�9�ORs?�1�.�u�RƸ���n΄��W�`��|.��kw���f$3#������mE
lh��`tu�%�8��9Z�k8��t��sV��+Qڊw�8�Χn'3l��6��9�aˋv��1�G�����ZS���=0�������^�����I�4f�$�<'���|t�FD����bG +Ǿ{΀�R�
�:9h���d�t�o����X~c3B4Y�WH7�Ӂ��P۫ �9����Zsc9e��Ҳ�Lk��w�8�I��{�r�7�.;s�'����"��GP+�3!�%�X�U{��S�&�4�Y}WE�O-p�����?Ǆ��u�%���1u�]Y%Mmw��k���c1��Jt��s(62ez��YHg�*f̣yM9�b�*RU>M%�m�ט/��T.*M�1��,�PMf�?iq�����^ܧ�B/�V�H.W�0�CimW�����\��� n
[ߗ�ч����˕6�1a��K�čk��f �������F��zYu&��t���W@9=�*��Tv:7�]��D����̏�
oELK�&K]���`�"6���i��})Z� C۞�Խ�e���@+�u�k@�7�[�t��w�1��K/G=}����9����^b	{J��4�����r���	=D���i�ŕ_�6شϴ��Q�H\S����F|㝟�æ:�޹�Z8t6��͙j���OwAfY\��]��FJ�j*�F� �@"�S� /*Ǡ-Z�N��_���^�`,X��[_�  �K��Q�}��l��XW)����a✕i�b���2\��Hr�fK(N�-�Z�����s��B�� �0��>-�yI��:��)"c<藛��:kg�	z��}������8;|�l���H}r��oFƓ�24���I�3ND^��]g��s�]H��D�Ns^��GA|-��툾D��E��#ڻƄ�#2}���S6}�e����_.$���r�8R�%<-�]��@y�A��UZK�0�|7���cf���x��'�X�ّ����X̒��y$WdDs����K[ϱ�*�U�i_�#~��Cx�Xx΁�u�|�