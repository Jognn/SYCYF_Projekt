��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&��n?��1ů��> K�-� �&�T�Ek/ֆ�\�놭5�DꢘP���+L+X�4��J��#�0�8���������l��jT��+�(���������6�MC!D�;�m�퓊D@v_p��䙋ⲝ��C_�6�Ռ��#�� ���	RD�4D��畓7���vn�H���0���fX����4 �CS�C`{��;�L����li��� y+����FD�p"��]���y��R��K�({� .؜M�������	^5���ɋ��&���&�@*���
e�� �t+���
_6��O<��7f�M��u���m(MrN����z�jL���@T`��M3��c�uQ�Y���%�dD���,�~^���y@Ga��(����C����	��G�86�S$��ɳT�ز8���:r��/y�[ݦڍ#A�����i�&<nU��<[5)�Z�-Ĭv���0t���d���"_���:�'-��d��*��q����_d�y�N-��~";#��������Y��؆���	6ZJnԷW��έ$Y�K�?�4���L�w�Wmiɶ��Y�?jx#*�i���F�m�E����O6T>]i�_�9;�!(��kH7�OS��_��[-M�((��lO�s�$�g�x7`��ZV�E���F��,9�j	@���]}<�ahb5~ãdl&I^�	v����-�@�@���	��!��d��`j[Q��� r��;f�i�.�m+UH7��/OV��c��������l��i��M��*'��?���G� SK�M��H?�ç��q;��)��Rȩ�"@���r��Ml>8!�S��L��EgeH]�8��>]GR=&���C��i�Za�z�,�F��h�q��^���wT�a���%�9�n��?~SИſ~�mu�OlIv�4'sT���/a��^��9��*��G�Fh�DM�_��CN�<�_Pg��O5��}s�%��m�o߫R���X�Q?��dK�Z|:�=��y�P�)�㿴��Z���^����ۑ�Y�t9�� T��l�G���^Q�F?W
0q���Xf:���k�ώ��H�1��/-8I��0���@=����g��[�;�vq-�%���FRN-���2�>Ӎ�[����S�Y� �ʅ��rHw
��d���۬���C��%��?��ES>-�|�5���r%�-�ٜ�_�r��T�$��a ����1I�kU�SKf���BX/�5�v&�=rx��`��j���ϵ�	I�I����=\�B ��B�M�UlP	0A����lj1��b�L���㞍i�!��Y�ݯ�:#�����&�ʒ9P*����j�W�b�h�M��Z��fT��]%���9r�}J�rh`[<i�P�f�/��5����+-�##���E_+&��3�.
�&9�f�r)YHJ�<l�&%��r��ǉ��\iaD��w(Xk�7�<Y[ ����[��X�>Yl=v2�j�M��U���T�@�����~(�Q[�x��&{�l.�&#0���f(GF�����qҫ��P}py��r�H��˫�"�|�95�.n��r`i�*G�¼*��Z����
�Y3f3<�ɼ���J��'&��`8�ٞ�|lu��g�ܬ���U��G�U ��=`�[���v������:�ŋ]���,���E>�T��lѽ�&�gnM]`��P忣�v���nc�Zj
f���ʩb���>B� �\-NXx�+z���qj�	������ =~�R�8�܃�`���*��WlR+<t'��(~\ҭ7�Ճ��bz �W��3�\�?D�\r�$��#6Ą�3k�Q���$a)k(ե�N���R�V��Sj����]�g?�E;��ɤK������l4�A�� �7f2 ���\n��#m1ɒg����K7GB�+ZqADE��J4I��&@'O��U�}(�D�J����n"4�>��A	{0�U��k'�B����N~�
�����2�b0B�%=>�㬯j�p0����Q��l�c�����YS���k �gH�k�v3���$Rr����u����{�<�	*��xA(�t�S?�(~�K{^�5[(F���p|%�����Ȗ� �"���.�m��j��j��,˟�[��%���V�� �~ɨ>�X�����T6����:O�:��_�4)(�T�t�}��{ϟ�28<�N���n
��X�?�W�J�c�o�?����0!���6bN6���܌v��p@kn�h9�ژ'/�D�Sr��z��`�6+wޣ?�Ȳ��a����%ȥ�!��hƯ��^N�l&������0�,�<J�@��/��!�5OA�}^瞤_O����|���KO"�&Na`�F��~7	�m��R�֟��o_�'��d Ή]҉y��M��I��h��S6}�D:��-����ثx<��fݹx����_x�[�Ê��Ѥ+yA�Ǖe��pz���E�!ԇ���������)i��Nׯ�u�� �c?T�?�W6Z_ï�ʲ��sq�r�#�k� �C �/o��l���P�k�[��uYF���%z�h�.8p��Gq�P)3��*�u��[f���D�MZrW ���h�}�2�VX(�f�����'t;V�$66�%�]�$5�^��/7:�K�b �R��58)&�Υ{�s��c׭�-�gw#�]���)�����6RvZm�R1�5���'��WG��l\0�f�~�o�g����f����%^C��5w��g��I�d�*�x���h4B|�U��f��'9?OF��8�E���L<3< ��gD����)���1P�
ÄD��$<D}����ޠ�D�����ԛ�9��i�:��O��F@���8��3�����K|3=7�3���)f�%J�-�C�g�A2����W5��8+��d�Τ�<Ub���ر�UX�p��ؑɃ���&���6]}џ�Q�L���Q��1�����$��������>U���k0�uu�l��T05���[��anL�~����$��\�ʉ~�j�U��=eV�kwBS�$A:��#(=����[��K��j����Pӯffa������{�]t}��@K�¿���@��MG�ʙ0:�S�5H�v�E}2	���c]�m��ͽ,�Z�n�:!�B}$�g5
#�ŭ��ȼ}���������o��I����2&�<%�!k��	C䶙�k��(���#�J�b���v�Ɏ:��gs)3&�~�/�X�.����D橳ub����؈T�J�S�-`���8�NN�Oy�ӯw"$����W%l���7З��α:�Wb �%�x���kw�Ya���g)m���@X�y�".���GF%��AK/�Uq��}]+ �?�9Ky�&�#tN�����[��D�}�8(��?�E
�㡠�7�T�Љ" V,�")��T���,��JK�Bq���U�KZI�b�|HU�t�r�+�.�Q�`�������7���� �<KVq"��`	�<��֕�L؋��ӣb�-&�����2eSl��2��H��rx���Z�}�g>�G+A枉����7���fSL��ŖJ�xEE36���~������j���HVl�k��v�#���&��O9eB��/�I|�&���^I��pU�W��<�1��Q�Վ:)�Y��e�k�[[3ЭW�MCm�.���e��'U������!���P�P�0]��:�|cC�g�03���T��J���,5��������H�k���ʛ��=\py�L.W64����koA�0w�˹ծux����Fl?u�MV~ag��'�q�8�� ��z��T�!iƺl@y�L�5���RJO�����t��L��26g����K�@�e'��!�ub�u-��� o/�S�AH4��R��"d�?յ�M��z0�j������;��x����6����=h�ll��N\�5��|�� �����]++(�NJY̓1���!�%�I$zt�~a����2��2�,�6�d�;1T�][��p��)�S�2��κ��}�6	D���� ���ե��Za���H�C�-7&'�\�"{&�#�U�vLO�iR6�� �u&��y��L����<g�V-�s��0��FJ�(�̂�����3ǿ��5�97�z8D�:�ȥ�_�9Ȉ�r���w>T`Òq/I�hp{S١,��zR>��G!D_� /]�?\�E�~E��p�44�)���z��6�����aO��s~~>\"��ps�7c����+@�v��{�qqyj�lW����:Lw���˚	،��-E���^[ZŬ��5H�*���A��<zǝ]��u�,�����p��P�Y��z]Vˈ��8�/�W<����T�����bmSґ:��*�'V��(ӒO���F�KRP�C�h�;Zq��<~z[R}����dsZ�6B����h��}J;0TÁ��x,6x�J��	������=�r9!�u�K�`���)�2d�T�ĭ�>��e2�(O�O��W+��Xs�GW�?⠷(��T\���}[���}�X���~H��#�'�V*�G��������	�:g��si�:* {�n�� &��
��n�R�JUS�O� �sb�GyR�Տd�yZi���Q?���������
�"�0�4�z��(+ T>y8�\xo+���i�L��P���I���3tR��iT�ߝoy�{,ߎ)�wj9�h��>b�'�i3��D8�Z8@oqG�O��N:�M��=ɒ��&Z�g�����?�+�9G��4����zf� ���P�c�@��'鬇�;'s�&X3]����u�'=��Ee�ڻ�N쎘k��6�Y�����Q�lb����O�����뾊x��2�tGc��n~㴌�ͩJ���o��y_k�Q��b@�g?����<���:P:�.�M=�RH�UC��O��:�r�����!F��G@Ƀ6�H$.R�����m{ՙ�cx9ɀ��!�K_��U�����a�"��k��˛���ǳ�|���F�8� �.����%�gQ.�"Ք�A/��� @e�b!��8#h'6�c}�-��2�!��n{<��Fz�S�L�C���M��N|�+C*�+^[T2�/H���q �SU<j�/�Q���>@uϷ�W&�i�.!?�.,Z�Q���F��C�J���5��Qhܟ@�;�Y�D��sq �e9���^7��>�u&q�Â�b �c��LcS�D� �A<Π��&�5��N-v�fiF��.z�R��k&����+�	��Έ�6�څ�go3�xM|����0����k%$��BK��+u���2�R��Z����I���m���0��Ѧ��a{��4QvZ��o�[��HQ����=V���-�Z��	n!�@w�\y�+�Re�{��	tm���~h�_B%t_a��4�� b��t�`G�|�YR��hwNF	8�uFvT�JO�=�*��6d�F�R��<KR���8�Mw]�˲W��P��q�͕�#�K��7�~
l��J��HuM���:x��Q���G3ӥo�^C�Z"@_f��{���r���c�����p>m����r���x�p��X�\cd�-i�\��F��M�}k�zOS�#��Bկ�}'� ���W��Y�K<�AD�C��YTW�x� k	Q06/�A�����hƻ��Q�J+����v���az6�p��#&"�J��H����mL�c^����H>A$K���6t�5�[?4��s��Z�y����`j{2�5
�sr ��"�*@��%�$�j?��<<�9�)��N�򗮚��Q���_ 15�L�(MQ��`]����r�J3s����]]+����p�A�D���ֵq��}���x�N�8n
7dAΤ��/�w�X�G�D�h4�!�f�6<n�����S��r���<%:-��L6`l��~��_��b����h�)ʇ����c����詵�3�q�Rfb1]���C��":Dk$<���E/�q�^+O�����E� ���M�ׄ�y�J,u!�d}��"B!��)jB�2ry>Y*V�������5^�����J�TJ� �<��)�;H��5!��.�a�Y}ѯ��������֞D�b���s���dZb�oT���H$�[ȏ�V��8Z��^ ����j��c���Ο({�N�<a��kUla5їv�|=� �uq�� v
~���.$G��ګ�0Oq�dS�V⊐%^Šb/��3�k��y����QY��͋�1���V�`P��R�A����{nõ�N*f�p��M
�L]��:�{��(gLg�ŋm�=p�-J�Dg^i+�r��z2�~����y�>��1��U����z��"�S��[P?ط�	�k42����g"J`�x�o~�r�����2�=�J�dQ�z�4JsƾPLS��������W�6�#[��ehi
Ǩ:U��W�'�0��^�O���*�E�Qfwl{��r*D޸��$}�܉�&X�*��o.U���/ő�a��BA���G)n��h�D	{�ڥ�(� �7a������6�/�;!���;�x���-!u�%G��>Y|gS��՟J���U���7H���p4�U��7V�yO?��#Q᳅Y{�������v;-n�R)T�o��{N���.�ߥ������+�Q%�7�]��%`q
���O��u��t���a��&�U�e�t&�#�A��,S�`�o�sgB.fU�{{{e����hӏ�v��HG���"<�F���KB�5�y� 80�\޸�Ʒ ͈ձ%kL�V$�b�[��k3�>4P�����%z�u���3��4}2O��-׏joF湥��V�`M�&���r�y�a��3�y�h9U�6;8g`�>��f�?�d@K`��Ra�����i�'ME��D=��\GI��;ݺ�����}�T>/xǆi�R� ��%�����U�)ǚĂݙG��D)���6gu��4�EmX�e��g{�DމI��T��r�U���MY2� �h�|ʲ|�f-���ަ"�f�U��F~�)N��5��������w-V�4���~.���L�.��b���N�����f�,됀`��l� 3��^�2t��Y�&��%2+e����� *zB�3(�����0U�/GJm�]8�L�
���.ה̫�+W� K�}C#ȸϑ D��LK�`��j��t@3f�v3)����
����љ�d���{��>�X���/"D��p�cX/�6/)�!"����Lj�[�!2�V�N�G��=S�f9E��{h�j�67��is$��G&۵�T��A��-R��]\��V�� �DB�[�S���%]F�-<H`\"��.b�Ք�|&��h�h��u^�7+�9��!=���v�SXh�x��5�u=/(h4��>\@6P��E yb^W���;;!��m�w��]431�nq\u�0S&I�����v��J�I0�=��T����������߮y����
m�CZe�ggH'���uuB�z�HZ�3H�h�o���<�e�`a���RX��[i�O��U��b�^Z�/�p����Uƅ��&{����=0T�e)��32E�
5���=ɾ֛�$ʶP�����)��mc�u��Ƒr�S`���;�?�S�edJ�Z�sZ�mN�>Iq�1<�Q������sE&�H�ٟ��KC�ei�����������z��qS�}_Bȉb�8��Y��9Й"9W�"�aU��AI Es!�w0���l�,�qd8�y;E����k)�#g��<��z\?����iM�`��2�Ϲ�����:vi�2�p�/;r�vz;�W4��Gd�ɶ�ott�3���V>�$����dp���$
$���!�����g��Btb�At��F��A�u�������<Ϧt �,[�+��� Ћ6o[r��F��֞���hV��u�~�t�	�Eʔ�%�S������t��R���Ea���4�λ�H��i>�������v�|��aO2���e��S�s��?����6;%�U�>s������YWk>/��>��@7�+omJ����p�(�ګ$-(�~U����Q��M,D
�\����B���]�����ih�Z�.l��o�|��O��%�1��B��g�kC�m2��/�޾�
0���+� 4����*�K->_)GZ���=�ހ1-�k�d�X�ʄԏ�/�D[-��l�i���l|]���3��"����M�Ƨ�ow�L��C�]�c�ِ��h�\A�HlLKb�:h��1�]�ZF�� 
�O�"nť���Z��i	au�����L	�n����Y��B?~�%�bh�U�ۅqB�َ��f��M��������$l2m�I��*ߕ�C��(�FC&�|C]�++
�^����'�M�r�ӖC�0��7�˶'�´`�C�ׇ��K�3��łA:�5�2��Jx��E���5kQ��)����u��"�)f��X�O���3��j���P�r)�����z)u
�n����l˜�(";4�� fF��ۋ�*�*���EZ��+�P�X����b�R�����R=���@ص1+�45����;,y���ڞ�wVe�vz�=�%�Xl�^�OEq��i�}$�cf�i��I<����a�k<Wք�A�,��s�Yb�?i����v�n�M4$G:��AVG��wUY{����B;�y���9�wc��(�EZ	ď�'F�/�������-��.2���L�V��]�ɣi�����UW�W��@�ܺX�U��g�b�z�'Bb�%zVx�ms�γ�1b�l?�}�I�2��q�W�qʍ�Wt`m�����7���5�q���c��R�L�ӊ~�Y�qS�E�R��X]2�}�VU|���i��_/��rB�"��F�TI�M����w�KȀ) �d��}'�Fnf��u(h]��+��f_z����o�2*�貘��š��0�#�f¬��k"O@X��m�r�(j_�$��w|�;g�X.��r��j���1�7{ϼ*�Q�R��*�ԋ/����<#>8`��wћ%�C�aRЁUk�����8�OOoY��mR?C@9�mt�!�G�*�� o�_8Ǩl���B��{� �s��[t�������'/9�{J����>��2P���q�SS
?we�W8]J�,?�^�2�N���f�Z�����m��=�V$R�@$�������@2y��y �>A	����Ear��s�r�MR�T��G����צZ�;�D��}���OAb�%q�!���J�9�a�GX�1M�H�[�3K^��� qn�#��G ״�˯\��o���l�i�k*g���>��Q��"���"��-o����}�[��KμMY�胎W���S�r�ٳ5x����al���?�Κv<���<�)n~�J���/�9��G����X��Ҍ�;���c�o��*��uǐ֝����Sh��1��nq�a��#M6����Y��z�����t�e��p�%�Cy�f���e�㴦�x�ғ�t�Jd� _t[nr�Sd�ֵGZhec8ٰ�o�U�v�M��Y�cW�H5@_�L*���*�)tq��$�Z%��4O�����4�g�s����M�u���,{3{����-�x��?�������z�aI�a`Xw����@�둌Y��0�c�+@RmԲ݉��>vy����(�$OW�8^ܔ�nc��8|^Pp��$C�N���R]X9�#l�/�tD8!���"��򛉻;qgx�9����q+���s/\2pݬ��!�n�X���e�S XLC�RT�C��p1�r��0��s�g2&�(�B��78nJ ;lG��b�뜵�S�ES�RO`6x�T�s@�����!��i,����8Y~^������>r��X=��Ɋ�6h���A�H*�r�<��t�QM����ˊ�^���d��2���Rv�zs$�t(�l����],x���@��Y��9�-�qYC[��(���tVt_$ʏ/ \�c�mMԸ%8�����V�>*ѳ�1@�\�d�s�ȱ�"`��Q����v��H�F����Zjqy�����k\��)I�����O������y�ШVs���N`�j }�n�}PC=Άs� ��|�e�F2��q0����`�Tm���8E�����D�3���h��ba�&K�R�{^�5Z�Y@n������E,�tL��|�e#����C'�
<0�qM�{ќ��%J�[Կɍ��� �������!���'������DchZ\�R�j���'D^��D1G�*X�����A�w�V�$��k���&̋ڰ>!����H�~�]���(��6e�O��v�TL�+I�:�+�l[%��}e�ۨ;MW�{o��B�]Wl��z���b�����^!G'ǈ�Yć��E��kGw���Ӷ���Q�N'�B"�����ǥ�?��/K(u���}�!jM�cO�H�óy��֦VI�m�
� �Z�@{)1����ЃQ����T��=b�<3z��3	%�6����]��W�oYx���[4�q�PWDcF�B��Xݞ��p��ѓ"1/���2l2����Q�n.��H�}�Xa\�c�v�}�j�c4�ڏ����`o�%yN\hz8G�h�L����W/E���d�]���q�Â�CA�{��&ǋ���R���eZ���H�C�!p�:�ԎBXy��B0��%�����8S�6��O.Q�ۛA(ua��V��P�s2J����+ٮ��'�In�=~�n�0����$�GQ�j;Ç�2L9f�ǉ�[O�&��0:(S�b`[y�`fRp�&�e)6zX��db"Rj�55/-[�J��$^�e�T�Y��o�&�wV(����?�RI��@�wQ�U9zX�q��x�J
b�ͨ9'��㑑�QMo�E�����'����t��z��kO�H�g�1;��7�W	b��ʋ�A��|�#�h�A"�÷+ s��u3 ��4���@3��I�S��%<�"���vX`'PJcu�
E�#2\_�(:��+�"~����)��_[%&{
�ċ.}��^��|�ߚg�H(�܉
��A���2�bge��N���y8;���#�G��=��/�R>��mx�Ō����M튑��ҝ�FJ�� ?s���>*��}�4K�[�1��p����6(�)�����)��/$��q�0�ԇ����w�V�F�*�1: ��FE�%{< wD�h�O����m�����	�ͳ1�Hi�JN�Na�R�V��݅%2NggZ���Z����#�!��W�U�`�a�I�~�	�ԗJTAWR��F�q�G:MW.S�������:B�p�䨬�;�v@�zYj��o6,o�c����=�y�.��ê�������,q9��<g֪ÎPːmwȘL*IںF�J�PU����\8^�!�S'���z�-h��KQp>�����z�-$��i��f��ܶ�]�pj�6����}�Ÿ��:rwc	���z���d�W��o����V�Ϲ�KP8���!�M���x�S�7H<[N'�b�'GḴ㟫č?ǑB�2����LĘx�{Q�c��4L�\KWƫ�NH��ɹ��p��c)70�6?�R��-��-��v�M�ۯ`�f�&v�
i�DJ'|����߰���ܖ���^1��ù��>���<����W�Ty�T�'EE^|��@�0܁�F�|\�!%DW���Wc�g�V ��mټ&��1�-m�Mm�[�S\>��׋�&; +j2K�,�Z=�N��7�.>�s߇|�ۛ��ƛ��m*�~�����Kf�!��)�`�����d=/��H�߷���,'�(���B+���tT�3�,�����<u���s���[���	=�8 D]a�T���B�j�R���3z"j9C�\85rF'� ���0s��2&k8�cUd���+M�F�9ڨ���W'It]
�(��c0O\E����;	4�$Z?�@t��&%�\��?�����Nc��_YغC7� �Jgʊ���|�L��Vf�C1l�kU�{����#���b���0��j��ɢB�:�6��u�n�gH��B3+�e��4���m�W�ܙ����}v�������3�_}���ENxWm%��V3�Zy~IY<Xv��_L�'��_�:GX-��ǲ+k��]5��W�>|�.�N,&���OnZ����A	1:<�N#h�f�����Iď|��у&�A�����������=��g���k�˥����3,M��G�\E�NQ5 @�=;lG���[[���,�����R"7�=o�X�G���h����>�#���j���rLFZ�K{bC�][��']p�{=̒�0��(j)��0��T�M�z�-Tf�p�O���"j �W�ȯp֡��C�z��xz�w�ao�����a��\O<H��@���Jn�玘no^�:�k0.�� x��OEe���.�WsG�  �Ϥ4Z�ַj��K�銽�4`�%f��Rf#
��E�S|j�`�l�[!��hc,�?r�sk�a�� J]�R��M�"XW��1�«��8><Q�`�m�C▇L�q����u#�[��r(_ò�d`�0�œiHV�Ϧ�B'��G<O)#P� ��,ƻ�(�7�<eVΰ���?m��\ʜ�.�����ٷ��OJ�0�+6`�3c�����Z��&e=IR�~Xd�P������c��t��>��Q����`6#�~~��"g�ґ|��aAsZ�]�j�n�a�!�n�B/�WB�S ��ˊ�f����i�r��4�SJ��f<
y�� �]0DD'�%�M�]���3�>z����*#���.�b״�Lg��Z[�k�� ��DX����XEc��d��l�����%F��|:�/Ӧ��>�"IB#���T���S��8����~E�x��Qd�(F627ꗜb���`k�fّ����b�<�߸��
��N���$%��Z-8C���pI�� \�p$c0I��M�ئ��mk��������i:�����Zc�F���ɨ�õ &�c��]���@9�?%�����7��攩�&�̧����S����i�޴��m��L:	k��浊� �h��5�q���-���Tc��i+��������sg)�]i�0��oӽ'��@ے�K'$�&Ώ�Y/��a	3�?lI��f&ZW>�8w+[v���M���e�Q*�mC�굦�m�YaT��g�d?<7� �C:5�;�M�@�Q�Z%�p�Ҁ���fO����w>��kM���u���LMa`Z�N�hB��}_l���c��.�� >	�9!�d'�&�8��S6��5�ߛ�j�vR�2�`� ��Ax��]'^�!�v���P��G���&��9HVs5�qV�qC����*�S������w)��h��EP�����\�j��N�����QANJKh�O��u ���[�0[�a (�q�����K�+<anq��\���(Sv��ne(. �
���O"��լmDl/���Q�wc�/Q��󥕶z�ZI}-�ZB7b���I)Y�A:qK !Ӽ$�E�\�gR,*��Z��>�`'��g`+�g���:0&��w�����L����?*]~:Gr:�te�& �����;�Y�ز���v?���x��#h���_���V���(���| (?OԺ�[��<\Z��w�I��1�����Oŉ��q�@:^�5�|K����)��=m*i�>U!���^�U['���J���Bjm
�ȓ+N#� ����fl����)��b��fp��M"6�x��1�mYb�J5����^m=6��m�R�NK� �e�[|:ll��S^mw)�	�C�=7.����d�Z�T�J������Kj;b�<��2��J�6��WX:?];	�ϲ g��E��`������\��NI{ ��M�)Ʀ>�W�bS��"�ȩ�\"���3�N\��r�5I��&벐OehRk�2�{��ߞ���{���T��(:��\�D/|���C��a��UpxV"���4��EI
=*_��El��j�t�`��Ӝ�A�v����#AY!���"q2� U]ead��}¥#YHB��
>;^Mmd����˖�;�nr�ub��_�0���g��M5F�J}����vb���iʒ��w��t�$l+�[Wϊ`����/ܵw�=�ri�V�«��U~�Jp_���5�bg�`n�9.!VO�"��P�GF&��ͺ#���Te�
������K\������u��>&F݉905��'��TW
b�����v�\��A0l��)����?-'B����;�|#���NH��T��^dY%��+�h��QQ�b���8}�ͮĆ�utr��qݞ���^�� �l]�EbЀ+�u�IbQZV�����z�k���]�B�u�1el�~7n��[+@j��?�7�C�M&�P�[�s+5M���b���J�K�%��T��M�������lD���V�r�!�ࣗ
��-��n%���(ߤ���w�y��ۋ�?��>	�q��#�O�눍X�9�4(�e�]������� Qb��+9�jh�'&�bq��E�%}� M�T�W�����ͤ��*�c�VOZ�ƚ��g�m�ٍ��Ϟ���)=J|]�������2�����������ai0Gg��6�4ڠ����Ȟ�ć�㑏��V��\6�J{��d����<�RPn���wy�)�b��F����+�%~GT>E������x��.C��}T��@��eohR�*k�U���+���vk!H�����a�Oɐ��"�����vW�AԜ�~cj��"�7r��#�'q�H!K`h�8�񪱝aVc���jL{�6�ؠJ$(�i�h��[4<�⤌�=��{�O�A�[W�9���[@�7�xe�\i�rL�Yڇ�F��8ŭ�?�9��)��ο]��Ȃ�E�{����^ph�'O�%9�핮ݺ5��g�J�Z ��D'ܝ4��ŝܙ0�"i�9����o i����>6��Ը�.�9�{!�¦FT(�X0���
�ϻ�d�B��ֽ�n$vZ��8�G���J�;
ڙ�h��»��#�8�֠���B�t��Y5,ƋO������ccˍA>�6��}�d�L��>c�j7sH��צ���U*B�xY#�m���3�N4�fM+�^����@Wf�޸�Ɛ ,�eZ�$�d!)=O�c�����������	#�.�\�Zb�����[ �O��et��;Kw�m�����;κD�WsE�9�t���Gq������_��0ɋ�I����%���$=s��%�_|A�]:�YL�����p.�G�0����@�C� #R��z[��0���8�"e=�h���(#����x�("3�'n�+lax�xD�M»-����@�}�J�;*���:p��d��K�$h���ȯ/[$��n�~?J�n��������s�3e�\����WeS��Z�a�I4��(�F��ֈ�@���m�Vr��㨱ӏ��c�D͗�O��V�T�ՈVf+�z��X�k��ÁG$||M�2?��]�[�Ii�`mS���$���9=��rv,��6�O(��gK+��w�y��3��X�>gӍc 8h�-���a������,:P�.�Z���7$��fa�z-���h�2K~����� ^˫�S! ���P�^�l%�<��-�~x͘p�|���|��Mk���8fAV�5k%x!A'<�>�&��m��s��<@H���=R΢��+��>��j
6΁�?t 7��ǳ07C�MKg\�Lzs�lm��|���t	�XE-��ن�R��@>�JG��i�'��M���yTG)t�Ryj�
(���c�͐�@���=�.O�xQ���R�i�E�8٥��;��*��iH�:�)��x��cV0s)�Ŗ���p�ߴ>t���Ӭ��7-(�n�>��%?,�a2��A�8Y�c����Z��%��;�UG4��r�t��[��#��ꆤ�ͤ�:�եk�5�t2
�u�����av�{
�8��MV:رD�lӨ���si�]uM�R�H?-O}��i�_���ͺ��l��Eu�z�T�7c{�!�V�s��&C�R���SO[����Y�amt�4O̶�L9�b�k��,�e��v7�߾��AW�%��7��]`��C̭8 ԏUO*�A4_j�1|��N�K��Yz�e%w��8����i�'��nh�����+>��1�<���3/�.c��@��l�=�8Ԋ͟S�J�9@Tԝ��6�Q�Y4$$��ZDz��mtuKR_��O���a�-�����$"�	Cd���U� `���'�aǓu�&2V�QOBy�Ґ�����cK�����{������!�J}�T�L!@�ҝ���� �{�͂���(D�%�(>J_�Ә~�y~��$U3�ذ6�[��1!�ӿj�+��wf�G�{*S1˯�B$���	w��a5qh]O�9'#������R�3���F�4�[G.���9����*�7�����]�@���S�*��j�=9c}^I�w9	��x����1[<`Sΐ���T!�v���W�
���%	bȮdD.�{���>;�.�5�4���fcT�����{6��.��qI�����s�v�vp�]kTli5��,4M�H�P�ʵEi�S� (d��b߄ǙsA�}��n#B�d��)���]�p��պ��c�W���g�͓+��s��Kl}�͖B�M���β�����-[ݳ�60P��-��'V�U��uA�
k/�4�'e�^a�U�&�"`��Y�x�u�L>Ö��)nܜ�ƌ�?P��k�u����W�b0�d��8)�R���8������*���`�ǉrʄj�˖DL$�w�9w��,��]��GF���%t2mЕ��$�BS<�1tـ��M_�*��k���!���s���&�5_0��J��/g����c���U���F�;I%J���E�M�ӳW#��mԇ�L;�[\ѢM�Ѫ�'mƭ3�V�����_~��8��5�H���m�:J�3`�zK��F6�o�d�@��S��O�K�l�Xĵ꿥4�n�Ud�W�āׅ���|�Gɮ�xE�k-|�\4Y�u�������g�"W%�LA���m�W?�m�L%`霉���8!���/Cʇ��q�t���*����]`La�@HPؚ�"~��1}��z8�\��ܶ�^��$�F2��u~R�*uz���^�UI��K�
�����I�X�i�ĭ�WQ��RSNVY/ZZ�a��}Ļc��Ph�=�Nk� <��2<�e��#��p!�YSC����T��I��U�5�+1��q~�sn��� �q�}&<���*��G;�Q����k��b����B�E���;JL�Y``����X����i�aR�cׅN�t��q6��e���jPs��r�آ��F`�A,o	q��ݺ8����;��X,z����|�|o>/��������3��~�W��3uf=���7A��淪n5x��& ����,o����57�Zϣ�ӟmf&.�S�[��l��`A�=d����ܷ�.�|���̛Ĭgfm_$���!L�]R
��*س�ǱM��$��5�� @Z0R��wD}>\P<�3�K[�D���܉���W����R����~V�����-^TJ, �����cn��YK����c3���f��)+i��<nI`��w���Y���%��^M���c� �G�|��tc� ��B'=������Da��?~``���>-���3R�_�$��Z$G�(M����D�	��r�b�����b�leBIW�$����dy��H�~ŷv��~⚯�/Y��s܁���-�F�*�B<n�Dz�;pK�� �k'�?D �\��U3� �h<�h�J����G��9]`Q5߳|�7��9#�N��'W�k4�,�G�d��y����QS
�#�4xv'M<k?��,��i0%�ݟ��A
��.P�u�J�X�,�1mW&ܰ`=���0�ٍ��A��O96��R�e1�䌕��[]V�M\"k=!�}M���2�F>��s�b�)���eY�gR�Vc&r�q��
%5���(��C�`�|��&�`jg�U+b[�,Ԝ�y�FYib��ut	I�x��|�)D�.Uu�"1|�r�`��P�⚓���W6�F^&���k� j�i�pgV�vL`V<��Y /nŽ���@a���5�ֽ{X#�v˿E���C���8:`^C�:������i/!����ϸE9�#e��-:���(���]n�g+9���6<��?|q�d6PQo�^�o�cM�o�E.�ZR;bC�i�/�V"�*����#MZHl�F2R�U�&�!,eq�=Ee�r:�HUwA���Z6��QDlR�s�=��J:8��-��h��� x�@��p�.�(�
jpUo������@�L�a���с���Ps���?D�5�/OM��5J��L����U�ZVWv�N`��h�w�-#��&�4�^�f��;K�TR�q��C0,���i|V�����6t�6�=*Mi����d?�P�wM�eO�
>H�B�:����_�ۋ�z�cp�"�^�f�]�7��Y�ڄ  ݄Xa3ɻ�W+K�Q~_RF�gi��D������$4��}��c��c�5" ;��T���k��Mw���9I.������3�?NG����� A����Jǲ��ޮ9�kg2A���Q,r��47Μ��^"	\� �ٓ0@؅j7G�F�ċ�=��W)C8���h*����gk�a9��r-33��_���}1����\���9����笂Λ���0�J����ȵ(�po��绮��Y�B�\IDw0���Ѩ:]�?��y����5��i�Kvr�s���Y�b��<
��{Գϔ��j���kb?�^|���]E�;�VdP֞t��>�	w��*=ggq �f����9��� x!Rp@Ω�93Z��)U��m���K8����IAcJ��+Z?2I����Eq���+|�jQ�
Z��	�t٢q���8n�E��,���#�������
�ج^�?���eS!�� U$��Oo
��@��@�~��Ț@�6���ق,�r��ZWj� e���ok] ���2tF/���p�;�A�]�;���@}/m(7��U�O^�(�C�2��$Q�e�A�ԘE��$�qX�Ư��W��T!�A�P��i�C��ȟ�v�2��D�'���Y�&�9�1̂SEbD�2��'�\,�� ��)����h�$�Ա��I�gصi��-r�YH0es�I�*Jo�Ai��v�I6!�J��i��/�Z�Z_�d�\d�m���mD�/p;����l�}����e�T.�k9���.�[�M��|�(c�KeXo �Hn��J�Q�Q�"�S^�h�����j�
{���&&k�NO��c�.��Et-P�Q�I(g|�%�[R���Qy]���z�Ws�'���`�N3[!�h�VN0�{O�F�f�D7v��0�[���c���-�DP����X��4Q��	�� ��nn��֏Ʊ�7=b�1����O�ߖ��!g���`�	�n9��a��Z��r�iqy(P'���ٶt)���W8�f�g�F�p~(]""��$�+8�*FȰ�z�W�e3"01Z�w_H�
~kjfr�l濖oud�N�!�fB^�UL3;%�����'�D$���J�*QDA}�Ɠ�>��h����Hu8n��zM�*������a[[������ލ\�x}דI�4��P4me��P�
�M�I�ON�o�]wUH<�x,���8��+�쀠WT��*Py�4��?/A߬n�uCo�n�bE�����c�e+��GYƼ,�� 4g���8l��oL�� ���@�6��{�n��S�k�ڿiSxOk��S�&�U2*�|�ieA���$Փ�O�Ǌ��F�@�`bo�*�qZ��6�,u�n��m��A�,�*�_�D�[\�?�~��e�����ѵ;߱uJ�e^�L��O@@}���q�gER/o@�B��R�-jb��?3���v%`�,w'%%0˯k�$���e��CAj�~םл��F� �j!e::1�o�m�������᷀�y�����Q7�s��P���L�X��X�u¯{���i1m�T�1w|##
������D��/] �ۣ�
/`����6,�M(������n�p:/��?2E�|��`P��Tb,���ȭ�e}�O��N�*aA�ˎ�a�7h�-�y��
�˿�_P'-�����!���3G���ܙ�|�d�_��X���P��AP���.�R�}��#@I��R���.�#b�R)�SBۨn����T��-|�i�'�(-�#�aB�QT�$-��_�I9�klJ(oʹ���$��I��}�4�~e�T�'��iF� 1C+e	�Y��M�eȲ�^z��4�қ(i�b���2�\�[�������0��_��ZLyo��^��l0����Ƃ���]�@�Z����W!���(=ΓH�
���:&��I驶�a�M��޳*_��C��m���BB�Y^O�&��7y�@G��D��1&~m�b[[�)��Gփ�@t�od�{����x����ؑ#�o�Z��7��8�S���W����0�w笭{a^�f.h䇫�l�kG2H���o�R��vӝO<9�Zh�x� ѝOi�ry�$���և�R�t2�{6U������w�M|r�&�y�3��)�a�Zv�w���
��65�`p�P/?�@��D&���oO��˞xm2����%X��B���j.�N=���9�2�t.t\�^��2�vwə+{N0>@+ehʣ�7��OQ�FA��E"[�����Z�R�ޖ�B�)v֊���6Vq��wr�&��5��+e�����M(6��*[��N���s��.��6iE)#d�;~��4��0�,�K_�
�{2�?��ǔ�=�Q��;�ːj�u�B�Ҫ0�3Y�c��� ;�
�^��	�l�v+$ ��#��V��-{����7����#Ҡ�EX>�"�SW���B�/!�㝣A��
{s�Q����z^��%?f��f#�fǿh@��1{n�T4OX*ƕ�u��U�F>�1=���rsjl�tHJN!�#Q��Ս�����Hm�E��b�z��	!Q��i톈tL;�*���i�-�-d��dlJ0�:�,V9,�������	N~�eTz����w�=��j��srųW�2Ҳ5��ry�O�>�-	S7l���o��8n����y�zF��g;L����C��]�V�N�-�Ey&�||�a�E��q�-# �u�#�+p~��)���c'� <d���e���l{^���]8�,�t(\W����X�hXm��H	��pNB>��?��M�U���q�!+HF
XbR�O���<�^��;K�a�I��i�%��"a4�ޖ��&���`�0{}r���$I������	m� ��)z�C�w#�������eQ�.ܽݹr��1]�MW����H��)S��pW�WBO�DL8. 9��&�sav�ޥَpH�㨮!^�)l{ATbZ�ɉ3�s��hϳRn_U��!MoL��d���`��l�K�]ȕ�?|*6�P��?|�pj������RC��N��A���Ͳ-#��̚���{�ŋ�PSG��D�]np�]@�ڠe�?ѐ�xK)��o�I0�ħ/*���h'���� j�����9��!x.�xvqYK���˗�<i�ʫ,5��j�� ���]
��a�5ao1e;�h��3l�q� �ҕ����u���1�;�54�}y�r&��Lʲ���#5��re-i<���D��w�{��������~�Xi�ݻ�ک�����~s�ކW����l}V)t��i�ũ�խ�3�I�� �x��Z���еu<8��}����<��*��9�_@�=3P��h>���1����$��^&,@(3!7�ۼ����g����°M(L�C>\�W��M�x�4PqP��.�ǞO�8��˟��0)G��/�� ��=�>��ڝK�4ɏw;N�y���>�*Q�|����ᖄ�,�f�J�5F�Cc�]�C쏖�vC��1�W�.{%t����I43
�]<2��ܘ�=�!����D�9��� �C������C}�죅�$���� �d�QL��9R����ys�#���ԝ��=�e�i�����?{ә`�M�'yf��
����7IW�@i��ב�&H��KӺ24Λ%�S���t��<ï�D`�v�Ї��i��_�-�t­���A��������N���Z�o��2g�\&j
>�:�;�6����黈�p�zv68��T�����55�Ɖ�ּ�p@0�j<����u��*ϕ����bX�(�E���Tg4����!NG"���9���rq�6%�B�i��ϲ����YN�c;3��t��yOS�.;�?x�a��7���}ӫ�3����S��áםP�wd�J"�uq�2�<!*���.�h�`!�p�=��{!?�cd�\!j���%�3��e¾�D"1[L�g3��n5��O�n�b�vPT��q��$�h��?�._
�h���0��������[��i�d�7�S�����L��b��������V�����H��{�<#������B�����BR=�ߖrB p��U'"s����$���5��̤_�^�kF�[u��,�;�S7D�}~�I� p� �>�S��0s!��P�b�w���׶�R��L�Jre�P-0���,P��9|�������xNK ���z\T�Ĳ���˄�A�y�D�^p�����#�ݡ��Ӯ��V�Z��mR*�	��=]v�-$������)8:�C�؟B����t`Y}�w`Y%�Q�I�����-,n�3�a����F��ND��zO͙�5���a#D�6�MB�7��r��$�-k+1ZY�J�XI=�rP�4�-7m�<�1<ItSU^���|(���+�6ZdGUL� ?4,<������'l/@PC>#��/������8��@�C���0�gx�xل�ea��(C|Y�} ��$-B�Hn(�ph�N�	Q��0B�褏x{לX�gy�VJ�s����&F��2�z#K�DM����R �������2��Ȇɨ",U.�b�c	NA����_�0��T	ĩ�p�0p�J��l��v��BN)�G�0�W� ���k�,��}���+KW1[F�C@��D��X�vM@=��k(]Wo��	ՋR�w���DP����2\Iӓ�_ƒp���~"��,���S˹;�IU �r ����"����G)�����v�AHT���޸�8~�G�S-
h��%e�͹��{AX�z�rv(��o�5ԗ�\0����8vS��t�3.#�]��徎w��n�������Y=|^{&}���f4�"���y:	$pSp�<|5��;r��X�J���|��������qF��=�����2=B��u>��QM�)3묵�9X��<#�O�M+�$�J]<�@H�ۗ8|����+�F��ț�¸P~:��78 ��O�F;A��!]|���ѹ�uJ	��5+�~����h��.�׷ٰ��5a?��UxY�}];���160&J94�D+4��>����1�Ȕ�x�$�����x�}?���ZGC�j����3~|�j��F�o0Մ'��Q!3OЇ���B�O�%w����r7Y��j䢤�2 ��L��n�	bX��	�r�N�j�M�:c��Sb�;��+lk=�Qda�`��5�&-�l��1ы��Ϧ��J#�X$�	�I�6��z�h�0бP��\kas5�hGr�[��Ld�*C=?�)PQ��ϋq�(���ԛ*|i���[@3�Z���L����}�0SH�-  =���w�;���1F�]���u�M��<��SY��cs�l�޿׃���~9��ŉG@xRR7�T���!�FC�3m_ON'���TOU���V�_��h�戨��C�0�R�S�u.�do��\"]��]�}��h�����pK�HO:�������rb��t/-u���Q5��oT����8$E���z��*^��P���������3隣i��~;�$����4����Af�nىn��gH����E��>���t��?d"�0;,���T�+\�f'b�+ۄ������ڍ�+]auUΉ�Y=�ƌKDQN/�3���t1���,C�;Ά�oXk�g�ϷזCD�V�Y mC�L�!S��ps@�����I�gc� ��u�c�u�i�����T���5}DB4W��`;��ˏ�?����]s%0�Q��̽�Xd�H]�.��к���A��s�1m����4i��Y�>��(���������r�tI�&<~�EHDL��B�������i�>U�<Zʆ�D�Um˸��5���_G����h���6��|e��$����مg�a��*&2�Ό�	�%x��p���|(�	_ӴM�K�4 )�7�3}��貟zm�p��ƶ��?-�l	�r��H���V�n�pw��E�	�>ĕz��y�*�輌t!�����!�_Zh��&��]h�(be��c����DQ�^C�]�U捾�?�>�>�S�acm�3Ekg��Y-���d���@�zq���Q��`6@��K9XP���#���۝F[5L˲�8�����b����Sl+��^�ǐ��'��P_��a�u�pB�x�'��SBm��0v�� e�0�F2���4������%X�QY�����};+ewF��[:�z2�vT�!�sii��H�������Q15�o�=cU�0�7�w�	�⺬�~�+��(*W�>��G��:t���3�_$Q��/�J@�=�$z��N�P� ߚdҖ�*��3p�~ 4Q��.Π�� ��=�aas�R���!��վ���٨��b��~3b�%-<���
h�Ӭ*8s�8�jY/#Y�:��!��A�`�G������i��F����"p'{8y��i�'�us��]�k=�G�ʚ�=n�b��D`�p��u&84H208�>�x���D(8�$ �B�����U$-_�&�豣�x��(���?�u�M��="�Jn��2D�WL��E�a��M�����j����4�d_W}l^��i�ɥ���ْ�=Y99�u_���*�H�� ���
����O�=ގ�n,G[ܖN�M�{k��o���jҎ���HV�k�P�׻�t�hD��8��ݴƋu��_K��9�Rj2�,��#�UQ�LZdS�0��A�pd\�����VHW�i `tfR���&*���.4��+����wr��'r��&�:z���p'�u�qۤ<��o��K�Y�~�U�3��/�UȌ�D���T�*�eV�����s�s4a�+d�Z�x��\�j�F�S3u3Ev�����5�.�<.\�r*����;n��%T�x���p�d��������d�ޜ���%;V6��������/�����*�u�)�jx.39�yX(Y|�l	{-ԑ�W}�ܓ�gH�b�\��u�J#��H��j�@�~֯"O\,�h���<!y�X��~���	���yJ8Z�{\���۞Ǌ��b���������=.���Q�2�V=;yQ����!e��<	�v>�T�N�9�'��J�r�$:��u�)�m��~���#�Z�e
�bz��u5���ݏI;�M�ȳVv��`a��Q����ļȈn`U��*��sց�g�Bh��I^�b3�{U2��y�6�Rؠ���c�Q�y�\�_�㵕�U���C�A�͍V7?�;�d�՘���q�P��!e8ϓ�w,�^�2�k܎$�!��Ε
��[t�����4�������Y~Y���S��G��`�@�� 1�k9����}c�R	x�Ls+P���Btvg�r/##~P�(�A���~2u�K"�	I����1D�mI@��.>v��]>]�P`�Fߴ;����gL���Ėz���������uX��j��2�J���c��k�f��I��x'�w@񢛾�Y$j�(�Dw�_9bT�z���k$e<ϓcjb�3�0����Rt���f(֪1V�E�?+�˿8�.��'�wU$+a�*���vw�p��%��#���]y�E��f�#nzK�2�j̯%��7��S˚:']_cXQ���]����擌����m�����J��`Vz�����}�#��=�X�A����.S/|���'�g��N#�_�B{��v�(b�v1��vR)f5:k�e�
x��o�{t�'1<�hn-�o��Z�8��a(&>��풹����a���iDY�c�� ��iQ#D�L��ƀ����h襒Ш�U���G�t���Џ���otTFF�bw�G��%��K��o� vn$���)�	��{0o@�H�$��t<��b@
E~&I���=�:J�����A���ǋ�}��pO{\�K���N��F�)��+���D��я&t�ސJ���'�^�B�_�
��R���ޤTRh>���G�9����d,Q���r���Ӄ���gyj��@q�ax �]	�Z���f屗ϐ��Jന ������z���֡�e��ˑ�����J>֓���8@�U$L}$��®ҿy�x򵹇�zcv���/6?�O�?t_Pi�h/4�pS�!��e��� ��j�UX���A@�:ނӏ�̸�E�k����r#���
��Q��Rp�	i�r
J"d)�h~����O���F!�B�L�������vG����	�`�KW�( 3���\��ծ*�\��6-
8��>c�,�qG{��4�X�B��޴^�c/��+���o�@��J�U���3�!Q��vB�y?xې��C�)^j��iY[c޵
Űy�<�V�8�/�k��� �<�z�Ã�9����v�˓yw �V�x��4U�ƈ���?5���e��^��=z(OG�Y>�j��XGG	g*�M��Fn���(�*+���=�Q�������2<UUYB���$1d����l&�0'���y�9�Уa;��O�Y��gO�����=ŃR
��Ji�@��¾ܠ�=!�F���`�T���/a�g��_���hcu<@�)rL��3f�n�K ߔ��O�B�W�7�Q�~�'<$�/>��woJ�R��Y3â����`ߑУ��h�OԦWa�`d��C�`�����8b�������@^�mͦYn��Ԅ�S�Է-6��Ra7��3�y,"j����y�Pގ�4C�ӝ�l��%�dbm��\~��}�����[��(R�i����ne� �:N�[����n�a�>: ���