��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&��n?��1ů��> K�-� �&�T�Ek/ֆ�\�놭5�DꢘP���+L+X�4��J��#�0�8���������l��jT��+�(���������6�MC!D�;�m�퓊D@v_p��䙋ⲝ��C_�6�Ռ��#�� ���	RD�4D��畓7���vn�H���0���fX����4 �CS�C`{��;�L����li��� y+����FD�p"��]���y��R��K�({� .؜M�������	^5���ɋ��&���&�@*���
e�� �t+���
_6��O<��7f�M��u���m(MrN����z�jL���@T`��M3��c�uQ�Y���%�dD���,�~^���y@Ga��(����C����	��G�86�S$��ɳT�ز8���:r��/y�[ݦڍ#A�����i�&<nU��<[5)�Z�-Ĭv���0t���d���"_���:�'-��d��*��q����_d�y�N-��~";#��������Y��؆���	6ZJnԷW��έ$Y�K�?�4���L�w�Wmiɶ��Y�?jx#*�i���F�m�E����O6T>]i�_�9;�!(��kH7�OS��_��[-M�((��lO�s�$�g�x7`��ZV�E���F��,9�j	@���]}<�ahb5~ãdl&I^�	v����-�@�@���	��!��d��`j[Q��� r��;f�i�.�m+UH7��/OV��c��������l��i��M��*'��?���G� SK�M��H?�ç��q;��)��Rȩ�"@���r��Ml>8!�S��L��EgeH]�8��>]GR=&���C��i�Za�z�,�F��h�q��^���wT�a���%�9�n��?~SИſ~�mu�OlIv�4'sT���/a��^��9��*��G�Fh�DM�_��CN�<�_Pg��O5��}s�%��m�o߫R���X�Q?��dK�Z|:�=��yw9����g�wd:�.��'M��<&6}D���9w"��e�1)-���!���C#2I�Yd������I��c���㭝<C�ō�`+UXx0����@�_M���t�L64�7��M�%t�X� =N�x< ������U��Ǉ)��G��24��>�7������P�G�F;�o�RN��� wi
�f����K{d��	P؁�:I�I�,D�n��QÝ��X���${�ݎb�_j;J*Fp�։\�.3u���t!mu�&�E�^�o2݆�������7e��l�b	���~��� ?����j��f-��3-i_��wZ�8T�ޠ�QW�#�TD�EIh6E񞺊�P�Č�m3h$�8�{Z��/i(��Ii~*��J=�Z)|�Ho��̱�PM�9]�e��k��۹�7\��"�[G�T�C�����\��k�,;�ri|�nW�"���
����Pr��`�oo����J�ᄦE��P�j��� X�I/�;0�8'��q�3��쾾��`�Xrfwvjx�#:�I���i��1Q2��]� dDVxph���ގ�����S�Q�>�5�ᰓ[K���Xk�6��+�� �������W�O�^�BV_E���:@9���3�.�����R.��D9.��˭7���#g�7����&�y�p�����u����H�������1�j�t7�AE��+po�r�)�Q�q+0�T-g��^�;D����e���}.�Au�����P���됵~՗�rS��En�Ѿ��L��]g���J��WW�n�6ŀ�������3!\L��lO�i��fOf�BoErᄅ4X��q���'y��#]����Yb#���ʚ{�F���4z̞��֢�����q=rQ<���~<=P�v�m����(}���_�)Vc�����yj����������76JL�!����J3�� `%>K���t7�1�m�H�f{���-:!N($__o���us��/-���8ț禪�w��몋Nu; �I��{v��l���"�Hkn+M������6�[��~���ݲ,s�Zk%��!_�������S�OU�kY��_����� m�9��r�i�<��*K!�&�1c5 z�u��Ց�< ;4s���D�Ռ=uB��B]t|G�hK=��Xƿ���_���L��_9�Qq[�_���$A�񼚘�K��Z/^I[�%���y�u'���>���my	-��_��e�uCI�i���lC"a/O��A'�>ǃ�{�W�#�|K��i�������d@f��M��iW� ?~^]T�s�+� �d���?��~�is�½WGZ\��j�����J�CN4������a�2;Lau���z�������P�%&'���T�N�l�?�'���6q�%r.:���g����	��>doS���^& O��O ��xf�3�k�]�Le�ȽZ��M�}ǽ�b�0�i� 83H��#���J�OrZF�����D��O3���>C��Š)�2(.�mF8�ɊSY����D_τ���|��O@���z�["U���
�6��u� ���D�5*V?c�S6�z�������2�� �U�tQhyY'�>q�<P�Z��ؚ,���lXɨ�}����U:�j��C���Nw��"S�K܊�(�<qu����}�d:��_-�I���ӖM��0����AX�Q���hP�+�$��,�5�8����M����++%kl�p�+���r�6��SPd?C�x���a�o?שUف.��ҳ�Q�� ��(��ot'aP�qJ1���X�4G:��ȋ7�1��������p���מ���>&�l��:�;,E(�J�����Oe�8����%�ޔ�6ޑᎏI��]�jG/iX����z���G���N�+8�Ǖ:��IU<����t�sW��T���_s��4k<��5�B�41�:%��T�0D�zm��咠��{]�q����L*d�b$U���lu�p��"cB��
�����^��S*n/�G��j[���gU*�rz��Ьo��^`��Y��r�����M#��6�'�ք����+>)��͜�PF��([�7O��=ǼK-���ر�`(cHzØ��[��w`աn(�j���/��Y�YV��M�+��/���+��i�+o����xk���?�^�6���ϛ��i�ygM)���Q�u�ϓ����{A�v�HoL8Z�מ�Z<�.%��M�}m�e#S���߷� �����Yko�ZOj�,)�����V�J��ap1I�9;��S�|��X�h<�ĵ1�Mok�Ƣq>	^Ⱥ����͜ ���<_�d��:�>ÑL^�j".$W%jQT ~���P���Í����u��n��QY$�uM��O�f;���e=��}��e��>s��Q.9y��ڗ(��ȯ6�\��g-�2_� �.�7��gs���n��L�;ZP@)p�I�4WHE���d��d�F��ۍ�S�f	��5�H�4p�Hx�[h��^ľ�?�d]��߼G�Ə΅��,5`W9|i���r�4Z<�NA�Ǻ����N���uR̾��e��ϹX^G�V��er�d������#�kr��;�c��ЏPO�`p{ �7�>'�[��!e�-$�]���	��>\��㭌���NJ4Is��f�ͫ�d��	����q�.���~�(���*F�N��[�nՎ$��H�3�Q�6���?�5=9��BNt�DN03�'J �+E�oe@�T[(.VEǆ�RH��k<$\�nV�E%��9���R������J!�%)��ho�Ze]��J�l����dwwᡢ�;bn��'E�s�G�ᭈ�|�Ⱦp+�ZJ�҆���U��o* ��f�k�9(9e���}�fhF���ݰ �=�7������|�9r_>I�t�����t�4
R5C�q�*{Ζ��T�p�/����5����5��j���hb	�6���rȈ�p�=��b�nP��p%Ŗ�V�IY��������e�mH/�&VXl ���토��|SN��Z���4��b�堐�Aihb ��Y��##7�G��h�м�N.S�G��GȲW��y�OPkW@�3��7O
��M�w�G�{�WO^26���>�ȯ�v��7�tL_���$��gJ��{s��
]���� �!A�9�<���L�%��7�����n?P|t��r�,��,�C~=��D�w�ӯ�&+R���·���/��Ê(��T�Z��HQBpc�`�g0�"Ћ�WA<��ƚ�(�J�]K?(&o8l����P�