��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&��n?��1ů��> K�-� �&�T�Ek/ֆ�\�놭5�DꢘP���+L+X�4��J��#�0�8���������l��jT��+�(���������6�MC!D�;�m�퓊D@v_p��䙋ⲝ��C_�6�Ռ��#�� ���	RD�4D��畓7���vn�H���0���fX����4 �CS�C`{��;�L����li��� y+����FD�p"��]���y��R��K�({� .؜M�������	^5���ɋ��&���&�@*���
e�� �t+���
_6��O<��7f�M��u���m(MrN����z�jL���@T`��M3��c�uQ�Y���%�dD���,�~^���y@Ga��(����C����	��G�86�S$��ɳT�ز8���:r��/y�[ݦڍ#A�����i�&<nU��<[5)�Z�-Ĭv���0t���d���"_���:�'-��d��*��q����_d�y�N-��~";#��������Y��؆���	6ZJnԷW��έ$Y�K�?�4���L�w�Wmiɶ��Y�?jx#*�i���F�m�E����O6T>]i�_�9;�!(��kH7�OS��_��[-M�((��lO�s�$�g�x7`��ZV�E���F��,9�j	@���]}<�ahb5~ãdl&I^�	v����-�@�@���	��!��d��`j[Q��� r��;f�i�.�m+UH7��/OV��c��������l��i��M��*'��?���G� SKٜ¬'�Wx�R�4{�ŲFRe����v2�	��t; i�k	�7
U�<��������� � � 9�84eL�J��"H�/��[��3xwlD��L/���	S��o���/�m����������Y����(rwNQ�2�nOw��رۿv��
�!�ںUʌn��3<�o�a���w��`+9�Sё�x�OU��}I�W�e��v�a�E���I�>I}�$r�&@i�ϻ"��s��,4�ZF}ST�} �x����=δ���^HR��OV�-H�;�5�\}r1y�E��{&C.Q��{i�������)U���C>���䚔�@�|��5�q&�J�u�b[�\�[�]�6��7b�`�E�~9U99��X�6ĥ�A49�8�Z�|��Id����w���z��[>�*a��0��Ӳ'U*:l���� T�.��Z��2���ϴ̈́&����2�>d(��*�T�i9u��_����_Wf��zV�����W�p#��ݖG=�JZ��
f�j(m�W��;��/s���Z��֗:���b��g���c.���R�.���YC|D��	+"h,�Q  ����X9���J!�n�����WM��ѯ��E�OQ�����S����|��X�kC^	�n@���x>�I\9�Q{�"�K3$5���=�?��[���ACo�����]D�k�QkB�P̗&��M�"� p�ۚ1�=U�xa�䫥�SQ�6��ils�(x���`hy�P��������)E����LP*]�4��{�j��	�7K;���� ��(�zV�*��L`�Fl$/�8Ob?A9��QTI# %AK���d�:���[�tV�Rѻ>Bl�"��"/�ӛ�F�7Ƴ}.�b6Wޗ�N��{�Z���qC<��.�NZ^��jc+�+?�$�^���R�UB�i��f:G�,]Y��>ُ�Υc�J[.y�ԡ�(L��U��	��d�y9����r�_9;�ä�e��3��h���}�ܰ�x�?[��e��t<��-�V�*a�����e�[�%�8l�a�=怎ۑ�֡5�I��p��|ŀ��Q��m�h	�gC�5s0��73|b6n�~�����t �V��G4����k���P'�dS��O<3$I�Ɖ�C ����K�`��.���C���I�ے+vMSnN#�p
��ҜR��\���]ڄ�����(��Β�N�HLީu�@��Σ�ͦ9�jJ�7�@~��cBO��j��to�@+03^ܫSh�B� �?ֳ��FD�ޡ�u"gگ}���ϢE{w[�����$[D����D�ϕN��#đ;/YVe�4�oǣ����&�-���w5�\W��]k%X;�����A{3l�@��B�u�;�GN������؉�NJ��Mu]�����T�9 ���U���J����J��1X�I�A�)4_é��C�*���\���X��w�f�C�^?���Y�2B�ؾy9^��p}��!"V�+
#?���w��ʏ�	�`�:;\�R
���*87N�KW;�Q�"{7�O>��vY�Z�= �%�Lz��TD�X�'�uTo[�d�MͶSy���L��mo�H�Ŗsm+�k�Iĉ'�q͓�!��FW�9�e���?�p��68��_ߙL����?�a��S����lFK �&���%'�)�ƫ��̊ZK�3���LBLP��h����%���@\�v�4"���&>�-�Cf�(+&��|>]�Y<^�`Nu��,���}��M~�@g��d$��ڡ:��EF���5��eգ7.LLI�}��r��T;ʀ��T�e�8k7����腡�L�Z���Ɛ��I <�%X��#h��)[0�Dc�}�8�����p#+˞}���9lp��\�? @��*�.��1v��.R��:�P����W��3׾����/-� ����3�W&�J_�z\���-��f)o�-�n�a���;���MWkL*�}Y.m(K�1�Q�e�p�u�=�\��h��� id�r=�����R�e�\� 	�q�&���\L�C2"���EP}o�NR���E��[=K��@�	zl��ڕ0�^z��n�	w0���M�uT���ިah�R?�O�J䑧oX��0�!��q�O�Ƙ ��J��>"��������r#����/��YlȂ�`�Y���R�1%��>�	�_3�Z�,��Al��y
_ȣ�Ѝ[�^/��ݨ��,�%�;~��aʶ���#����tM�ya��Ry2�E�����<�C��O�5��];������w���$)~��WiF��H�'95�ܴz��w���;\�y �߯)�5�e�۔��B ��r-��
����k6?|_����-���	�U�|�l�ZB:����t��_{jV�Jyz��
��xF�"��JG]�V����|T�����*Z��F�����>'����Jpv�Gu*!����LY�ɡ�c�����R	a�
��?��ҽ2Wtۯ9�Q�8�����S����6��Um�^4��&B-l��p�#�"6�F�\����ӎ���!4��ް�^��e�|G�U)cL�Gxzk��oN������i�^#H����AYY��5IG(>�b�?2��3��,�� �ҵ}wxv�y��\�J�V@�6NG%��T����7����rQ9�>~l�ى��MǛ}G������?y0���l�#�XEux~Mj���k^�J>�έ�;���5s�^����r��K�l�$�3S`D�a`�܈5����3�n��H�&�/�t��1[�a��%'���p�[|U?��ȓ�2Xb�oi�p+�~��ez�"�v3�!��(�^��m�-I�2�@#%��e
�* ����j�
�Ǣ`˩�	�3�$y���U�]��9�<��s�2�PUzuu�;ʐ���F�t����N?�]G�A�"�xo�!y�O�T��
�4���t��y{	�f�2Fz^=4++�Ƙk���AR٩W���D�/`��>Q�#h[��L"9%��
Z��+���6BF;2�j�z�?�1p�wX��(&L_Y�@�i�U�wd��"�'�Flz�q6���$B�R�%�w�[yc��k�r+27K��t���~�ƕ<�ʜ�Ƥ�=����X���K
�oϳeP�q{�^ ���H���	�8�F0���c��G�3ʼ�������{��[q������$öu��Ϩ�3p�H���L�����=ڐ��R��5�dq�1d"l@m�b	)�C�̬�ھ���v�(�����u|�GK�f+���u^`u%�p�I��'?o���ц'���ج�����$ڸթ[�[7Y�^vv\����ʴ+�[5���L�q��oؗ��m��� �����♠^�R��D4�B�v�b�^�}�/�����3��i��{�Ֆ�utE((�}Ps��+�U<nf�?��}DB��`u;�P��^.U�8�kK������-.�����{��!H��:أd���W%Qy�kʏ!S�C��p��|g�s7���1�g���#ܷ�4F9lSNm�(���`�J��3,�{1�\vK�/�is�Η.h���' ��-�I}�_r���O��T��������a�� ��)+Iջt�Fա���]!�������0�.um���`�k��>WЂ��d�I�E:�Z
���aͫ�$T�@*�)}�n�@R�8]1	R����wP��`(�u.`��0�ô�R��2�]�W\�[S��d�� \hup+<2.��Hb�q�Gl�4�,k��A�D������=&�)����[�^�܀���mVb>�6kۨl�ν6$ٍ�+�q%�\�	_ݾ�2�'��M+T��������'�2ذ���+D0�.���p<�q�U��|e��@�θ�Ӆ����W=��u0�[�U�s#��f'aT��~���T��B��瑮o�Q�Џ.�-/ۖ���Ub�!Іs�n{_�9���!�V��/Z9��SX�C�5����p��Αi��K!"�o��0R����F��޶E���D[�L�Y*��R������5[6�P\�����~G��v�\t����|�j���=�� d��ܤS���Hb�(�>�L�����næ{�̝����/uό�,*��	�����$c��>ֿ������0��l��^To��Y�!�	�ZH���q����'��(�����j��P������(��^�;�	w9,��B'\I�*Wc���0o�D0Z�d��M+H���Z��gz�������� �_2����'>���Ţx��)�`�����X�$)���ҭ��o��z�)�c�
��[ Zi�fc�����b'`�ٹ��!�g��r��h	Z��p[e�MSo�ؤ�f��|\����9]��(u\�.. gM��K���_�W�UO�᧐������i�z�j�l�X����| 0�)�<NGB�8������<2�y_@[��h7Bk���n�Ww�^�-�!�ߗجj$��6��$���B�H�WC�$"�OH�����H}<��pK�N�,,_��J{�����0�WF����${0�RPr�p��P�t�F���z5h_���=��M��Gc�^�o�h�"��ϰ��z�mt5y�;.Qp>����U�]��U.2�7�o6{}�e�~s�������D�����ji�����Y��|�ي��~��z�o#ذ���N:X�P9Fނl~U<�����\⼸Rb|��Y{�����z���.Xf�KO�}��6=~��hkuW�|b!�JNs��X��@�Ď1i&�C�Ӎ�ݐ��Rc$������|<��)N>���>�9�ܴ�����>,]��!�rt�=t#F�J�O�~	b�DCF�v��l�Y9:6M����X�I[���fA>�v)Dh�t�
�y]���"NN#�T��3�k}�J���bg��!��xo��_�~���QD[n�K�1 �a6��S������}�����)�s����س�����Z�t�������v�O���z�v�ڲ(���E�ҎV����pz��%�k��s�2�[��E����i�I�C;�b��ux����f~��A�F��@��@�k��l��,v=2�ǫ���)(��P��Q���=�-N���񢂫Q�#|4k΂38��,̖Z�3V�yKC�h~F,��d�.�ap	FC-=0�����b/��k-�ȆyP;hbM[Q�9�1T����B7 ���x��ϑ��ۥ�.ƹH���"TMظ7�R�c��&&wM��baнn�]�1I��Xj��nӛ[���� ��+���u��p�~�䋓�����<u�zl�x����!<�(f׿�����vx�~3�u[\C�k�6D��ҝ�P��_#P���	�S(t�B�w���5�Pi|�V$ǒ�����v�!2��&�i�Jmv�nN2�-!��m����E+_��qZU+6�M,4����1�Y(,���S+��|^A�P@߳��Ϻ�:��#�ZT�B!g����'_�y"��h���X2�u(X��i�E߾暁.>r灓�l)���<Xћ��9��`�(�vZ�w)�s�β@CkȪ3-���68��b��5��O���F<=��S#�&"A�C�#�����DM&��yzl�5���f���C�j�^`x�X��iH�!��n�x {�x�1p}���2i9̓�����q�\Y�gR>I���k-�Ѭn_��6���D�Vŭ-jP���L�94�?���|"{�V��+C��Fl�j|cǲ��o[���b@��D��9��#�S�-�����i
DJ��i�P>�#� j�b��卢����uл1i����F��(.�y)pg�
�Ʝ���~T�{*ߨƣ#�/
��h��;��E����+���>�ϒ�����k�h"e1�&X��s��M$�6.����9?ݴX�ݏ+�3SeWM��X�Z.�%�,y��	������A�m��ط���s��O1�94E?u�%
K(�syɎ�ёه�% ��<�䪱�˥�W}&z�;Rcz��uo-�DX�9I��ĒH ��-����`=�`��^�M6h�u	�"�{��;�5�ueo�֍U��z�g��r�υ��mK@�X��5���ѯc�b��!�l����}]/�'�h��!�>�h���[��vcˢ�����~�p��?3) ԭV�	�e6\WQ�d����I������sh�8�.��P���Wƒ�zb{���*rIu�$���qSoj�_���i ���A���"�����B{3HT;\����VHZA�P6�L��ӺZ�X�!��)����kz�06 @xë�r��pe)J�y2c�S�>Y�.����蒶䋞d���uH)"�&ӇƜ�5�	ʴK#|L+�������,c��q8ȏ�S6�E�.
 �2)s�o�X$.�}hPR0MTe{�c��ҶO�LM�	.�J[��"�a�!�Ub�F���*���t�Ɯ?�{��N�64S���x m�;6�#��G�sM�?u��"��pO�F$��ɏ�i�2�X�AڣK�9\}��t'ƻ<�x�pw��oam4������K��O������zi^x������ک_�Ōk<���6	�H�MI�v.g�A��Hk�&C�r�'I (���։ۅ���V��j+뵇l�)5o�!+ܨ�9Tʏ15��$������⾉��vi�_3hw��Ih��C��L�;ǲ��"����
���_d�)@�Mv����%[���^��#��F~iwk�9�v���l&Z0�M%�/3�z��ʘz(
�&����}c�܁�=�{@E������<Yc���J��>�WF�>U�l.:9��j���X�?��4�>�ّ=S!ǃQvEY��(��P9����ߊX�^�v��R�>��[f�#~� ����YZ���IQ�*����A�nAcV�`ǖ�?sP��ػw�����u�)$;���E�AU�� s����Q��m듭梅ڢ��9 �h���It�t	�P\�Q`�?����/���gR)���xr�Ҧ (�E���?�@Ǹ{6��Ej������[���Ntc�T���yb=���x%y�>)-�p�l�o�K������ρ�(�O�r|N\���VX���r(�^c���X2��7�Af�u>�j�&c+�X�D�U��Pq9�?~K[%�w�~� <����}�<�M}��~}6���Pm�W s\��ת�p@Y� ����C̐��V���7������q��@��<@�e��Ѵ ���.W�l���9m��\G�?<�'���]�ZƜ(��Y�`#���*�@Dq���,��F#��p߱6�,C��21}Cr�,|�Ú7�ى�Po��wN$�XQ��g�P�D��N@��� �`�!�6(���x5saw��U@���cE!�̤+�q�%�>İ]8��Ƈqd��]s4�o)$�g�ؖ4]�غ|�����x���̡�G1Kc/
�!��*4j�)Z8�x��ϰ�ç֪�8v-�uM 9o�[��Ԉ-���!~��Q��_��D	��ؘ�);��mmQ-	���lbY4����iuXb�_�=/aCu�LYm�F�>��KeC�w�:-�5�=�3�KW�E�y�����2m��Z0��.fI2����S[%7֝���K�Q�.��g�;r��bO<LZ	��%o@h�w�D�-	B*��^�3þ���f�;
��[M����2�ա?�Yo!����i����YV�}��J�lt߽F�p�ҲF�c��zf�t��Kd锆����}�N��B��+Ix>d���Q�2�9�BbPW�9?��qd���������˄��o	�)ut=1H�}���y}�h�!"����$mr� �ds���3m�l�Fv��_��l�֝0����-��P�����p<�j w��'�'w�u�J�^&QY�d��W2Z�2a��-���"�G�<M��!��'\/4h�J����v��t.y�Z}^����̆UZ���lQp곉�Ӈ#�姣��
�"E<��5�æ�W�%9͈!�UP��a�B����o��H���S�h"	�(�	>T[�x����-�!Ҽ���c�ɑPęDn�5��v���I�˅�'g�ܞ|�7��� rЄI��f1v�'�#�
46&7�`��Enf2�>�_U%�1��^	�`�4k����0j�l�+CCxnt�?��!x�w����7%b�:���<g5�0�$�z�T���19K��0XZ�ppQ�����Zp�\.]FPY04 b���K��|�ɰF�Z�r�9ؒ����v-u$�E��Ҋ⾼���E�
����G��.%pIZ�v�4'�By��vuUU�X�DK��1��4,𲵆@�%���D�����7Rl�**_��:�&EAaA$���L�ܝ�����yM,��co���B��yh�?�G��>j)�"!��tߋm�Zr����h(�i�������K��.A6���i��8SޏS�����x�P5T�)x���s�G�7O:�B	�~<R.��ř{��w	Yc�:�����������MG�A?��}�#  	��������������g)������<�Ι�B�;�s��r�ވ�^��Խ˜��޽�:w>^�Ơ�V�V�2��������x�	��
O�q����u���}o#�D��a>��r���� �qW�!�����M���F- �BUeL{w�)+n����DGu�|�����EP�o�Y
a�ݯ9���p�c�˓���ǡ�aE;������P)��������'��(�U vّT�RU��|ћ��c(n��ϒ�W��R���mp+"�t�Y��S5�<���J �s����q�gƻn�l�k	D�K�$Ꝯ���S��y#����f�"��ʭ���б�SZ �Z��d���$�Z��W�0:C��Y�rM6lm|�)!+Ӟ����m�H�Ŕ��˼�W~����M�����Y�Ij�ڋe < �C�Y������%� �6�c�� ��X0Q�C�Ǣ���?��c��'*�RU�ヨ����@�܎��?�{A��V����!e���y���
ț%ݓ����`K�o@K�Ѯ��q�� /����Z�'#�����,�`�O�H�\�S���o���B�<�'Ķ��0(C��k|�q�������@\���ޑ���e۔�;~�� �B4��^g�GPo5z���7�b�߻{>�Tez7����@Kc.�n�e8�WRf9AG]{�����Ա̇�Q��w���NI6Z�kÊ\7��e��!��Kxp G��rh!*�-���,�gE0G!��U�'#oG�ʊhs�>��tx���]�3�l8�R�'f��&���;����v:ҿ���/���J  �<��n:%|�'V(p�vKZ� H˒4qaz@���9AB�K��G�~H�L6�d6o�L0�Hn�����Ju��HB���h���8�z�]��j�\�vٮ��Z}M�X;FB�Ȼ�<K�2�o�0'���2��٪\x@y�|��3lHp�-��&h'��L��v\�q0�E~]�ō��&`��1VL���U�ihҙ���쉱�sta�y�@����*��R$�H@��q�dc�0�"�o�O������	��u~�M���tF:9�K��pb�.�<0�B�cR�A�UXG�ܣn��s5�W�O��r�Ѥ�06�w�#_�<&�^����2��V�� #�B4' ?$��i1r�&�_�毭t) =��d��Tl-���c0������i�"`@kAc­-Q⮦�];�>.�^Q��j5k|t�/���Lh Vk#unF�4�f��_���� ��I���zḋ��چc��;���k�ڳt�ON�n�Ҩ�Z�oEo��������8>�?苽r�i�Pt@*p�|����&�����Ĺw���'�훽¿�^����2U�b��U*j5mL>��ÜC�X6Av�9�T��c�J�7�z(,C�_�z�����q��c@v�����s�\���;���#�=�L o(��I2J�Rȋ:*S+�1.�����-���(�3�T�~'��� u���	�C�]f!u�ۭG��?!����/6�k�e��TmT��S�1f��Ē!Z��Z+B�q媅5ï�W�$�������y��2�-�J����cWo����U��S&�~��A��ޡ���5G�Tis��ꡠ�N������{�m
G�� �ho�X�& �.�Q�{�W!�зQ'�T$�3���rPLn8׼�6�9�F�KgZ���NB�̀1�~�u���ۼ�����bp�wN���&nv�m��h���s[���Y(��z+�7���J���{E��'�����8��`ᚯs?�~G��#E�������C4A������/"Fy&�ڏ�6b@jS�#���6�c��˛�y�$�t=�YD^;BӨ�g~N���B(]��<[��|X�w@�o+<[���w�PE�ζ ��&���񇲌�J%y��i�k����;R�3�=~3���QBi�!G�r�ɾ�5�3�����Fݝ)��8����e깐r9�v���\�[3?��D���y��7)��4�b��D������+��S�# �;�������!��;7e����Mf��;��y����L��t��T�S�j�US��ػa�F�_Z%΁]�}��� Dcp_lq�VWD��v*8�h���cz�X����E��B��$���%b�9kͥ�a\���,�K�N#��[�r1nY�	C�����+܍a];`qZ��%3c�V���άE�K5��{� g��Cw�	
ʻ[��xH��{��=�f���9ZR�������g��)��
wu�gg0n��p�+��+x�!�E�Vwūv��h���"ːC609S���&y�o�Bk�X,�׼��,F�0j�G���Cd��u=�ʰ	�ҿ $!�T]DTP�����V8DA��E1L�w��|�R	�`��d�]����0%�w�,*���}���t9�fڋ��n�2���[i��v ����e��ŷյ��D�+T�m�ֈH���i���	��9�f��hu�?G����4T��)�,�B��n��+ �Z��9���匏�xC��� T������	��v�zs���݆��S����C�O!X�8`�)��"���s��� ��{���AK*1B�f"N���&�݌�������kP��n���?m�=������,�L�p,���,ى�1dEL{KIU�Qk��J�����Yd�>��I�+�%�R<���{~ꙟ���Y�
\|LF�.�ľu�1쟬>,�����<�$�h�*v��qM(m��R8��d�&)[�|�݀�aV��Y��+l�ɜ�R�}����h����Pk��"S	��j��kŏT��+��L���ߌRKU�-��-8��{�������P��}3���Ƭ��
�$��B��:�S1Z{�d%2�
ŭ�;�����u��������ӳ�c��N 
�:`�U��+r؞A��i���qԾ��(��c�4?�j�X��:����G�k%�u�28�(�e��A.X�:KEd��i]�3��zGS��))m�摣��A -@��d��ℐ̭�po-f˺�$�ٖ��9���'�:�r{��|�Ig��`I��3>\^���t�R�� S��l��h
!<I�����T���w	e�,�����Q���1n�2��TGtף=�v+,�E`5"s[�]:)$�xK x��-E2�˘b������y�:�f�To�~�pK�l�M�@��<N] I\�]J�]6e�,�w3N_�y�R/0����[�8t~�b�����ŏaG_��	OEy����;8_l�gD���dS1Ӊ�d)�\�M������m���#�r��F1��u}NVO3����p�|�&�{a8�gz�&����EfI�S fU��pA��hM;��L�K�a<w��yτL.���m�?{y}5�����ܸ�
�0�2�<�A�2<h	Pr_�@`0;V�hH��ȀP��b4qj�L=�T=��JvR�&Bd�����le_'\0�4���g���[�{�v��O��}��ҍ��@��Xb��m1�%a�`Z@�m�ֈ,�
�{Ҟ��}�
�<��Y�����O. �5�ޟI�(��x�y! r��uY^�×{�oT2�T�[�~[���rxؕ�Z8�xQi8�P��p��"��d���I� E��2��qd/-.�7gқ2�P���g^l����>V1�=@X�,]K'\�j]��ˍ��a_�|l�A�����	�Ú�0>&��>uX;����nfXo��;��#�٘����a9v?��.e-v�X%��҇�
ڎr J,��D��s�m�0 �qS�
,���C����43ff�XT����L4�Ø��~���l%��<2��ؿAq�3}�cM��=PE/���U+�3�b�>:���,��	�O9�V�TQ7pZo1��g��Q1�u���H	�(�:e�ʡ,�9Q��[s�IȆq�g��ވڕ�j~��͡li,'��41E�ۓ��'tl����ʅ�^hŜ��U���"��xa�y�I��s	�I�$4��f)�x�X��x���j6�@b�e���)�h�b2QH���a� �6��/
{֤#�SiB`�y�����~�@����Rro�)-�,CV����z2B���'�9���(&�(s�W`M�ܿ����k��ʲݓzM+\<���� �>�5\����dr��?�'�UKC���=38��F�b�@�ݕ��I���%;ҰD��w��u{L���J~��ޗ�Bd��~�}H!���&��q₮5�}�d�B�rI���ܣ�8o�bbC��#(<c�ht��a�y���]����'��f8E�
�@��&lM�=����Q�q�=[ �&��["�B��V�#��`������ZaכE�[�>�BS��p!H�����o�UxN:���OT���x�Y����չ�TkI����i}�Y�	�&���?��!:�с�ɿ�>��[����7D&Yf�����m&^�T���L �����Q	.]�����?�E� �]a��,��;���ۂ�>(��0� T<3��}�!ۧ��!��a�5k	ĭ@��H�@�*3_�-���iu�S}��yŹs�t��U~�q���&��)��1�+%7�IM�j�����!��u�۽y��z�	�F�]����"	��l��d�/���T8����B��MY[N��]^0�
#��W��<���І�Ւ�6���+���<�qxWF���]*!������}�9�­ч�/$��������p����h��rT�1ș��$�hP&���넣L�/Y;�5�HܽV2p�[3?�s���� yۍ��kՖ3��B)���U�B�c~	>K��5:�67��Ą-��RD��|a���+J�c��ھ̙��(�Z;N0N�QR|]+�~5E�D���� 1�`������|�c�s��Mmc����<ϡU9kX�_lI ���n�� ����,~ܤ�)�y�Y�.Ɏ��0V' n����k,%�Կ��4+j�ԣ�Ê@.�ܑ����b�������j���P7������&+À`�&�����0ܹ�4X9ل����.�D
7�`8jGD��ĥ�����s7���x�7������z*��%�uz���l�|�Vg�����כ�VQ4O�����1uuF���u~���X|�3%:�_��jB/�ɦ�%�Q��"Z+ߢ���q�F��e�TPYkr�Ysb!8�G��?�W8��l]FV��@^����R���J�Ӯi�oOQob5�`v��l��{��<N%G"�_�M��p^d������;�(s_c5�|$a����rv%��'բ�+���xP���(�ľ[�@����vYw_��PPB����@б����,>�G耠�#�$��D���<��mniK@��Ū��5�k ��ø��}�8Rx�ro��V�7re�Kx�H�?0~⛖�sXKg\�����FD�,��<��ܗo,E�6O;\��Ȱ��pS�^��r�!2�}3li[��h�"=M����]�
A!�F"]J�R�ⱨ��u�y@�u-&�/������cu�*7y�v/-�VXY��tۃ�C\9�A���ܕ�1B����S%B�L]6�JZ�ٛ*�s(׽��8Cf#�&B�.�u���}�8][+ Ln
��L�kf{�q��7�k\�.�JZ��L��T�Q��N�u�7�k��q�MM ��t'�M�Mh��+#��WD%�����z��T�{'�d8���d���K��􏃘�Oxۼ%^�鴝hU���S���r�l#8cJ��j�:w[�D�3?�r�n���Jᷢ�]y��b����T�b���k���Xh9���ra|L�T���l�� �j���3](�
����i%e2�:*ou�~�x�V�5W�~.=Q��e�{T����"�%4,y����9��V����o�k5޻_m��$lnb���T��k�T���Ġ_,��hĔe1�Y�h���I~�3�O(sD����/`V)U+�����Ͷ��hF������Vߧb��<��ڡF"�e9{��ƧLl��sZ���c|]�]l7��WG�BL!��3OG|˚@<���ǰf�S�5�64�|��h��ݰ)��o��r�;��☛0SC��
˾���fbؓ��>��M�l#�^Y���y�p��^fj����aR�f6Za9�~��Ѡ�]�A�V�����Gb��H�F�{�����՘����M��P�^�h.Ab����>�� ���S�QX�'DH�u����'��R�B+3�i��8�z��6vm��x;uF2p\���[�Tn��B�s'�4*�N�2�	��k�tJ,�L*V�kT	x
�������S��-��z/ |&؅��p}o�8���|���{0c�qQUv��I<4�.>oX�)ґ�T��X�2r�P?SP9s��;o�3|��8`���a���W-�6rժ�	��~���D���E� ���ou~�[/Ɵ������o�e;�ڬ�J����Ȣ�I�}�gl2�w����+��������L�Yv�B�_��w�����"*���R�R~T�yR� ��0��L �;Y�9[�� rY��'��X�\s�ԒN6��f��^�뢩��oԶY���,��x�T��ܽEL�4��a}��%ɪqF0���U�/��$�i厢v��*Dc�ۂ�FZ�TeC��Rx#9<����?�<�jl�P�AH�w�h�T��$� ����n��g\ܶ����?�2A��f�� ����ŶN::df)�(D��=Ϲ�$s�Jm�� ��ʜ���Ws.�j:Y[Z��"�|cB�l��C�Tt_��Z,����t���=���"���Gr��c<�"�Ɋ�B�u�E�$R?vm�ċ������|v��;N��#zAB\��_��:30���������X�Q���n�Ʊwݖ��I�~��m���Հ����fN2�S�U���o���"Vt쨟ȋM��%�\�I�_���=�t:��Q�~����6��0M�p0����Zd���Z�+�5��������%�g(��U�X^=�_2�%�R}�����\�g���Ұ�|���]�T�� �qPHN�U%�&��{���PT[��ڡ#�2e}�w�\�cc8������f�g1I�ƍ�A4��\�U�Ք��z�)k��I`#��^�L�]ͱT���|i�u,�c��-,�@N#:��O�dBs���2Y7Z0�X �t/_�+E�3� ��ۤ���HBK�ڪn�xJ���w��>�RA��֦z9��|��w�mp4#�������+���P�a���mu�;z(�Ɋ5��'�ؼ|r�m^���bX����X��}��� �h�{P�%U���5P�� �YP��`�)P�qE���%���w����gw7�Zvcg(��P��B�%���� �z���"�S��O�k�y�/�C)YxA�#�!9��q�?O/��L���[�}@�����7"a� {�q�aF��~���tlcUdb29��8�8�]0;���#� ���̀���j�>���^/���:������@#�WSx|Y��,��*��\q�OE�n�\h��Q��O+��kS״��q�7�A���z�� 9�ج�d�,�����䂝iϖ�29uZ�.0].L�5��\̔��O\��'��=���OJtt�#����yBk6U�\��9'�1��H!g�sW��"� ^u�:;��48�U$4�� n�7g�G�wQ����!�ij ���$:��S�KG�힇CqL�=V��"Ӌ�k"���[�<z�����1B
%�-��u��Od�H�@�|v��$�/O�cz��a����t�ٚl�c�M-����f��4(�+mI���!�-��Z٠ϼ��g�b��H�3�X	�ܯE9x�JR��8&g�O2�:�0[Íy�˔�!v�r}�!F�I^wd��������BַOn��v
��W�zq�p�ذ�A��w��zIDI�����O"���&�j[��o|��n}7#c��uK�q��O���a�Sp�Q��1�����7͞sy���2H~�-2�/Y.�h��d�����T���� J�&f[D��2���c�:�z �s��n���t�7i���:A��M߃V�>�S��W�l׸`��f�!��S��Ip\�XP3��x�r��N^�!��|�^�	�3}��h���7�L��h�bQשH�Q�.� ����Z����lxK�{�JU%Sר�L��Ʃ�v�[�RMx�+���&n!����q��E�$qI�Ppm�w�"�+J��W#���fU���P��|E���@��Yf��&z�����Y�H���Շ96v��^��(��ߛ)�E>R5�{�K��q/����Wb|E(E��+�y	�0�p��ۅ\N���O�>���9�O M��8�x�+���E������-Z���?_��q��I���R����Zͩ3u�&P��^���00���o;�6�')� ��]�����7��XV��\�tPHxO�TB��j�`%����3�/�L�����Ρ�p�U��2 �<� /���(y�E��D����%��[��9�ñY���Q}�a��1�#�QG�<����`�zX٥C�����R�U�CL��-F%.88��`��$�_�ikC�����ci ��O�a�×�>�_1dC�=��,ɮ��g6 ���`M��5󷼏����{��Ǯ<�H���~x�i�R�]_�(�k�G�_\��&�K;��j	`(ԝ�*������tD�rA����٪��W�σZ�ԩ���dme@"L4⏱����Cl�枴,Ih����?�p�虂"� �~~���έ��>�W�e�a����k��7o���|G|�k�#�[>�V�(����Ri���G4����!e��V�2>��ĲB��"�i�u�T��r����<���?6kr���f�*�N�Ǡ3t9EmVYc���#^$L�����=�a�
E9aÎH���KJŤ���*��ORU��:�	�����;�c�۽�GjH�A.��V��F܀��F�����a�n�@-i�ax-��7���,K�ﳹ?6/ԩ*�`	ey7gp�V'^K�������)��	�.����n����|Z�UP��v'�4��̭p��ɅL!�
�M��7}T��A'��QT����&^k�9�72f��U҉Vm�ܧ��
�������A�w���$����'�rB��n�r���Y���H�dz�d�<�y]�2����M� �0+�N,��I��Q�|��̫I9����s/��m;�ܶ�Tl�vЂ�!����QH!�>�:�y�C���OnH�3�K�H��� �f�x%8��Z�5>�@4R�'��w�a��-5s��=n&�����M���d����l�b������2k�D:���l_
!�$�^��r�*KV�m�Df*֪!��+iز�����Qj+>�ޝFj��<��w�<LʥU�h���� &�S���;��,� �O�nﵤb���7���gd��Iu�;#I��l!1��3�+p�~(����[IN˘�t����G�RsN�O�^vaY=?��"�����`���+U4�踪�]�M�;��F7H���u;{J
[l���Ӻa��/�
�r\�4��<
��Ql�:	�O�t�>Jn�M&����ۇ�\�C=[F�ء�_;���,١/<�VA�U{h��=@"�(<��
�8b�45!�j�u��C:�fiQ4��+N�]��;^�=J���LF��ݎ�7��U���>��Ž1AU�Zg��Y� S��9�	C��nLi�&�!WR/ؠ�QIJj@L������k�=����l�ގ�~��C5()����Ӯa����۽R]��v�����4�sb�"�ۡ������b�r��"��d�ðn�+�� ���Qm���b����`$�߶�m ��_�����6?{.�Ce*�x	d��i^�ٗ�T<�	L|�-��X	j���t�5��y���uL��:��)SI�w�u�ƙ�U��ݷ&�ࢄ+�� R�ҰZ���"gZ �b����Mq���i�^D��P�K�Y]����e+�I��P��}R�F�)��&���.�д[_(ɰ7I3�Ͽ�tΖ����Jj'��=��]j](��%9�-��⬀8�&`�nD�x!�r����ׇ��J����m�*rn�T5 ?��;��7�
o#�F-e1��z�"n{q�ġ[k^R�p�n��JIȥ0��|-@ع��q�������`�:Hz����!0mg�����|�y�?�])	�����j�;�a�2�#��F��D�U�,<>�ST�秺$u�)y�/�2��紶�T#��֚�y����1Z��8n�:ǘA�V�Q���E���L�
�4Ի���h�t�n�I�w�����˘c�}!�ê��|�	�,*��.KE�XK~fR��kJW<\� ���d�0�:���-����S$�?WG����<S��ʾE�~>���R#��qQ/�Y��h,��pܯ
��oՊ�g����E� X���G1�d�~W�y!����'�eQ��;7��B@bO��S�-��;l@�+@h�m�kj�s�?2*��G����*�e�Fv4�䗵ye.d��q�Õ��x;TD��W��D�R3�ͮ����4��^YW�lR�`]<V��rɍ:	h�p1��v$�}����*N��D)����4H� �� m�Jh�o��@�6�)�ȉ��FYƩ9+/7b+7����'L�zq�H��+�R��h���z#a�(�/�6-D�)0�#�?��eW���}\�"�ւ"9�'���x힏Tۯ��a�E[�w��X��4+r�;9|d����H}p��#VM`x]�m!p.c���7z�%7�#
�0gv��+5���L���wؗ�6囹�n<�@���ar�+�`�&��R������ L��	(ũ[5��וpz�*��8$br�՞�k���`�Ў05I"�T�c�N�0z���I����'�#�����:|����_��i�r M��>BN�@�l�pFT.�j��J�R�"�"�)�g,%�_<��Q \Ə{O���$�?
x�$1�}6�ޮ�����+��P릉�w|-}��JYX��bw��y7��TY�GS��̽#x�K�B�{̾<6p@@[�HR��}��1��ޟ:4a�b�k��$��?������f�8���*�U��Ê?�*�P�gg^�� \O�@~�'�$�ƫM�5�|�����M���M2�ų��a�.M���k�=�n,1��e�����aw��Ջ�Ejxmf�Ŗ;)j�����	�z�'y)/{.D�?�UX�e{2�~��u�8����)Um��c�W�N��r�d���<���J&�Uȡ`qB���/�^���y2,�	%��q��I��pN�����S�
rv�e�0�_�FwO�.�%)�y���g�R��6�.��B춸���SE�*H܁W��#����^��0���R�� ���hm+�2���@A�A���[�,�%/l0��@�A0w���6�&O����x0j$�f&{&;O��;���������N�w��q�4&`�JY�`���,|�F6ZeN�m;�i�x7���uky�L;W���:��#U�H���k(��fLZm���2�a}v�L���+����zd�UL�.	z���Z�w�.�rM�>,�����G����7��(N���]N����N��nBtm�9��ܣ�N %���(/��Y��|�� S��1�Y/��c�[E^�Ǭ0�\�2��?�FP�3�A��$��N��.1&��I"=�g$��$��*.ӛ>N�PO�G�P��q��笶T���K1=�y��8��G�2���6>��%'����[�Ϣ�|��h]��I۳�bT��q�*}n%;V�(�(��"�+yC%�!}e��=�=W�`Ee� ��'
��+%��I��t���v�փ�qQ]Q����"_?ޘ��>P����d%��ڦ#Y����<�V
����D��xg��ӵ���� Q(1�M��C� m�T!�5�D�I7�9�'�؈^�J�T���Gv��4�'tV���]}�)?�\�%s�A��>��������5�P�Ӭ{��ƓF�$-��$���)B��R�q�J,R���傰���Ae��'B�+[�X(��p�;���f2?%�v����N���d��ֽmA>rDqN����Ķ���"���ʭVoO����9����n�3��Kϓ�^����<�D��	���k������e{`���ѝg�q5�*;6g�Δ���Q�v�E��鵚��W+^�,AF7�-��*YH�*J�i��;2?K�q�*�s�W�͵����ɂ!�ē��NUX�G����_�Fk��k��D�yOZ#��K�7����nR@���i�Ckb���B�y1XFC��L!g	VK��0�ˁ��R��~Y���x��)�<�Q�)��-��Ҩ���\��z�.��29���l����D^�2���Ⱥ�c�k���>���QGΦ([��*nd4��!e�[�JM�$�H͏6���9��\L���A�ĝ��b8�_Sx`|�,�鬣q�V��
�I��4��B.Z�['F���̡�"\ Qɢ�ϵ�JK�����m���S2�*������Z��b͡)[U�c��*"��2J�����%���o�5]�L�f���)C;��Vݠ^�>Y_�ǟ/[t���>��&�H� ���9��'L}8r��l�1�{/����3=;����v9bn�_�Q���e_�Dqf���m�����_c��$R�"֮���	E��|�E�d�����"k�Nt~�BI R%Ǝu% w�@��o���h,蚡���m-R�a�]VB�@���>F`�}���m��M�4����2V�Z�����u�A�������l�]{氨q�Gʜ~��5I�R�7A�!�ʾ��	,x=7�C���2�'���Oʜ����nO2Y�Ds k֬��u�����v.$�<P?�x 	;U�
cH�q�ug�$:ݥ��a|��HA��Q���HǅkaS����Ø��Ii�^�7z�od�`���Dd�ݛ�o��|�:bB�[%�kԂ��zb�i�-�Wu�}u_�^��-�fk�g|�و�Y賿A/_�4��ŽѸiXs��0w��'�6�*�V����kI�M�݌��"􂘑��(v���7c�x��9�&n �}�*�oe��0[�M -^l�K��P��@#���BMtw ��,$��b�ӣ}p	�wc��s�E%�-�6�;�Ec�����?�ڃ��o>K|���	�X{lKc�2���?���Mb�5���:H�kR����0��CO�9��F��R<j�G�U����o�W頏N ����6��y��X����π��Ć5�S(��������.?�Ǳ�hݒ ���	r�R�
�7�B�p�?�D,�Tq�݊�4���!ұl�q�������>���K^�/�*z��&�G��.?�ٙ���f����W���\�XPQR��F�G^1 ��8�ܠ[>�t&d�Dn�Wb$��rgȡ��?b�Ӈ8{E��P�m%�c�z�"�b��j1Z~�x����9�?������I�L��NͦG��m5���#�_����o8��/y��޾-�`