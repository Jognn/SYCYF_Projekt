��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&��n?��1ů��> K�-� �&�T�Ek/ֆ�\�놭5�DꢘP���+L+X�4��J��#�0�8���������l��jT��+�(���������6�MC!D�;�m�퓊D@v_p��䙋ⲝ��C_�6�Ռ��#�� ���	RD�4D��畓7���vn�H���0���fX����4 �CS�C`{��;�L����li��� y+����FD�p"��]���y��R��K�({� .؜M�������	^5���ɋ��&���&�@*���
e�� �t+���
_6��O<��7f�M��u���m(MrN����z�jL���@T`��M3��c�uQ�Y���%�dD���,�~^���y@Ga��(����C����	��G�86�S$��ɳT�ز8���:r��/y�[ݦڍ#A�����i�&<nU��<[5)�Z�-Ĭv���0t���d���"_���:�'-��d��*��q����_d�y�N-��~";#��������Y��؆���	6ZJnԷW��έ$Y�K�?�4���L�w�Wmiɶ��Y�?jx#*�i���F�m�E����O6T>]i�_�9;�!(��kH7�OS��_��[-M�((��lO�s�$�g�x7`��ZV�E���F��,9�j	@���]}<�ahb5~ãdl&I^�	v����-�@�@���	��!��d��`j[Q��� r��;f�i�.�m+UH7��/OV��c��������l��i��M��*'��?���G� SK�M��H?�ç��q;��)��Rȩ�"@���r��Ml>8!�S��L��EgeH]�8��>]GR=&���C��i�Za�z�,�F��h�q��^���wT�a���%�9�n��?~SИſ~�mu�OlIv�4'sT���/a��^��9��*��G�Fh�DM�_��CN�<�_Pg��O5��}s�%��m�o߫R���X�Q?��dK�Z|:�=��y2�}�.瑷���}�^
z��}X��W�>��O�eX����N�H( �]��礅��O��U:0��6;9�Xkw�O��ƻ=�*~p6���	�r�+���R�6s�6�)��O���k��y�|��0��T��Z����7�@�����\��4�Q���Qc��3��ٓ,��YrvX�w�A�N���-�K��+bh/��;�SA6�cw?������.�.JY��h�)m��ݥ|�'�,����X@7�"��sm�F(����{�r��1��[��dQp�����X�iFr\��Z�� �ռ��D��qh�4��tA׳��"�S+dѪ�*ä�c��i�Ž���L	{Gր2���n�R�`��ݮL�����ze���\F����Ц Ցܑ��I*��%I���|��
���UO�
�X�y��ڜ���;��)���-��Ð/�d��P��CxS�-o2y��F�~6�V���:��I�݉r������!4��dS"�j7�����,s���/�J�U����!'��8Hc��V��]H�#���7r^��~�z�#�$+:����;M<e��0������Nt2�^{�����zc
��}l���g��Y����m`&A�4�u8��r.�����3b�[�k;~qb5����X��
����d���&�N�lZ��e�Ё���	�ֆ�p@����R�/�i;_{��l���n�o)^�(���ڔ�f��9FFZ���m��n���
�'��˧;(8	��[(d�B�}5�=�] p>���+ً�̦=};N!�`ӂɨ2�'��0'ݗ�O&>뾟q3���v�d=Wx�=���t������߈[���y���+(�}��7Dŗǂ��i�﯄Z���#>���>�H��H��tp�xV�`���(Z�A��?]^�����A|�.�ط��xg��Gxe��P��?�p�A��.��D��M	�k��� �AVUk�̺`�g�S"XiZ�wD�>�h�a\����nMԢ�������'�DPJ�	ڗ�"<�ž$n-fF�K��V�zKmˡ=4S�����G��c�:�yU��AF�i��"2x8���6�T{&W���3x�$��RU ������&�UG��B �R�$�	}X� ��v��a�2Ԣ�F�ɬ	mt4m{�M��w���L��A-F?��x���HL���ϙ̮b�����!K�M,�[%�����ߋĨ���ku�
���p)��r����c*�ޙ�*|}�R�xV���|���h�O��@�8���#����#]�\�4H�|�� ��Vfԟ}l�	��r���0�@JQ�!�YyC;=+�|��; ��#�
Ч�@rܰ�-��΄�F�Ƚ�G�����@\��$�w��6z̍�� ���վ|���6e72W���.)R���Ebsp����I��rb���x�iX��Ty��9��*�r�;��Ȥ����Y��@��!�C¯��h<�Qj��������x�Q��iNcLw���*�[�<�A���"i��G��qU�o��+]Wk3���p?��l|�]���0C~)s	�{�,;>ur�;�a��~�y_7�7�h�suϻ;��^��L�9���qΎ��;�!�6�@�'���t�e���ݰ��7�EM�ے��?\W��f�OP[�'���I��ǈ�G�У3�9H��#޺���1�5ء��^D���b�MƓ"���=��GD��Ö%nc��s@q�����w(�}����P�*��<������y��v>��bAؾ�7��(B�[���%�h����E����a�T.��P�r�܍�j3�-j(���5����=��@'��9QQ�i%����
�g������&�����>�Gv���:�Q9ޙ2� ~�O���/˒�/iu�RԝK�E���.�9��,K<�)(�1���*l��z� 4��Pg��}<Sd=�?]r�"@��׳��~�Uʲ�O4�Y��9��ƂN]՜Ȩ��6&�f)�����;��,�t�GB����&=��F~�#o��f��Zx茕�5} L؅����੒�l#��3����l!l��P�{������m�X�b�-_�fɊ�#/Ks�x6b`�}}o�C�an&V���#С�{��L����TF"O����_),i?A⸭��˺�?F_����4vg�H&ux$|k�R�N�$�iK�1���G7:�{�EǄ$���+QD�r�y�Z0���.��:�C�+�5�k�mX-�y7Q�/��&0�D_�;@'���j�#��1p	�j��^�MS6�,��#:ſ�~�ic&Ρg��"������(��/�W�y�h���{�f�@ �G2f���� ��v*)j��
����>ՙ�q'g����7�9�@w�9�_T�%E��i1-�}��2q��>��\t���6��]c	P����͎o U�����~m%�ɛ�SKM/l�bb�����&�	�����C]����u���0��`��L賩�� �yۥ�+j����ߋR� �.����$}�o1�AȪoI���{�}�A��$�d2�֘4=So��+�z��s�D�!r�}&3�p���4o��z�A���^�ݗ��uS���t���-��4�T����d�D�TS�X�@ Q�Չ��]���d�ƾ��Ε\r�H?�&�G�}G�⪠I�m��r�ү�B�'-�V��q�ب�Ķ�Z$�.��5�K��O���y[���
X�a�wҲ�Ń.��h?��e@w�\�����AZ��6R���FaNdAߎE;;GQ��J�8�u��*�w�u���9�oCMo�Vل���m4�ަ���BZ�1���e��ޟ�A��S���� `?b�6jsU9��kG~��(J��x�Ϸ\���`���)^��p��Wr'(E��d���e�s��y�G�����n��N*�/�iV���-�"'�\�?�mK�ڀ�Jęf;����
��L`�4O�T��ˋ�;J֞�b�Y����6X!��y����7�"�KQ��'���-��\��a���,�<��4Y5;a�ϬD�X���+H�f��nwfp���MaL���[��+��t�%!f
̣H� ��?�="T�z�au��?v��-�I3+c�~�뷗�S��l��E��Y�C����08 �Ybg���0��d0�����?= q���OP�p��L��<�����d��[����6h�Z�|w?j���ݡU��r.�hM��n�e��2���[ѡDgg'�q#���)G0��i.�,|�ڌ{֏��;}�ß��B%y]�σC�b�O
)8˞��?u�_�]8|ϋR`���������ߞ����n�w��٧���ɕX(
�U��������d�.l���"Ë��#KQ6x�v��s��;�@�P��(�a?�6P b��J)�J�"f5@l8�[��R��WB?qs�@��c���p�<��3j5b�����t}�U���
�e��m1�bFCzX~Gz��"0Hr�FM\��֑1���$�����}�k�������3K�T�[Z7@SF%%n�_�|�Q@j򕅨���M�\B�$Z<Wh9�U+�ix��}��w��pK�za�*�P��͚�J��G����J-}g�f,�h$�c;5���K��w��)�G�W�ÑSڛ�⛘��8#�N=�K�g��P�k�8FNG��!dƬg'c�JD� ��j�uN%y�(��C�[z�Cd��W_8�[mN�Χ-�� ���a��Ե_��R5M�P�5"�~jثQ����(Y��)3�a��T����ᰦoP�����#_�Rz�O���5����M<�b�-��;��~���15�X�-H����朔dӯ���0�cv����N�TnI�Sy�uo;�S*��aaS��6u	4��y`�OI��S$Z�Bs��|���/�:XB9o7�'_�s�3#<9�,�EO��o�������#ڑ��MB�Xp�
U'}��mD)t�B�8aIT�(��S@;v�`�:7Li6����~Mȩ5����e�p�����������Y�K" �R޳�d2 ҨT��*�|�DR�1����/�
�|�/CY��o�$�<`=2���'���ը�����g�H�)t�ek^��!��� �!��9��f7���y�u㦽S��J��<�v�s�4���p�(�q�4mR�z�0:��5z�'� �l�>R'���i�y=���U�"ǽ�� �c�N��=[.X�+������w^"�����
�q`S�)^��Apr�B��m�f�Oud��G�Di�p�/��QQ~�/ũ�Q�pXr��f���r��O�x��|�n�t��щ�d��|Fi^�~��!�U�H�j�\Z��70�zwP��ZT+,r�D��3������=&(*��c�yj(��]�HC� ��ڀs���֖h�3!�f����@D��d�;�r0i�!"����E���|�u��9��a[���MOc�Pˬx�� Xu��L��U�S�2�}+U�ï&lL`�`67�/�wOϊE;V]v�e4�]00�*	�:�KYw�~b`���|��ucj�^�Υ��T.����T����I�8��QB|��AZ���B0"��b%��ѺQ@mu��75��C���l���O�����s��/Y������1�d��~��/�e:ʗ��CT�c�$va��u���IM4��-��q�N{b�	��f�IU��pi��cB�2S=�5�Y�H��:*oX�ʩn�efo층Yǩ��w-lP�BM%3�cea8�Y�|b/��q��*��k~�dȯ`���w)�� ⁇QX�(M�ݧ��VO�!�6Lp��q{
��<�a7kD��'��Mqi�ъwK�T�@��R�I�k�,��+ҵe!*|L�:[9'U"㥴� ���Ӑ��s�<³�p��|�~�	��|=�d�P(����;O��dWJY��Z=恩u��L��0�$��:3���NU��	j�ga�Ҍ�VԠ%y���]�K��8�#�~���:����ħ-�`5h9no؊��ϥ��	ܑ?.ۢ�i�>�@��^޸1�BH�x�Ok�{�����4�ʈ��q�R������͔[^(���w,�ߕ${������΃����Ƕ^8���$.K�C���,ع�(�d�)��६�u��9��������#u�C0�b��v��+�"���נi�p�L��}Z��Eo# X�cv�}�xW��N�"��-�(MY�D* ���}}Ƚ��v��򟷉�7�|7'q����l^PZ���jFы�4�|��[�kv�䌳���
�@x��a�>W˕T�Qu��@%�1K��	D���#�����>�� Q�1�X��޽-�zǫO�����}�/B�?&�rv(�byih������ƺI ���ѬD�7�ux`G50��|×Y����gc^��S���PLJ~$�J�p@~<�+(�X���,xt=Y�O^��0�a�? ��Y�E*����s%l@���m�)G���� O��RP�!�B� �ìov��H�Z� n��kc���	\ֶ������}?*v~��26G���9���^"��uVT��r�cq1s�3�3�L�m��A<J��U�����W� *�W��ąL��čYf��ɨs�R��x�Wc�al_G����4���9�q���M�oTE	cc�Q�фN
�0p�m��´�b�A ���=ч��ƙ����c�@R����b�XB���wW'gp�H�Xb�@�:��C��.�X��@f�L�ɶ��o�����<���ΧLP�������<y��\IW\[�O��J5���A��
�B�2���#5��G�Uf���w7�Jr��%��%}5qB���6��)��[*�����䍠���3�Z gׇ��2�7�ښ�kh@VK��c�Y�
w Yh�������5�Y�
;D���޺�y���UXX��WtxO�v��kF.ÂZ�4�[�Y� 8�Yhw3��^Q
8��c�Z)��B�����@t��[0�6� �ݳ�X0fc@"u:J�D$WX:��*(+J:YC�$���~%�[���� Q����[�:Y��m�8%S��Fg-"E\���mg�{�1b�O�Ή�����cw�E�QI�����-a4lb�Jrx�BEQ?�`{):2�Z'�\�c����n��&]ܶx#{��&��$}�n�� ��MIX�Y�|�0���5V��	�}}�8��*a~����\�	���Ep�{*��p��ğ��d$'�2{��ne^W=]=eW��<ɧ��1P���(b{����r��Pet�G;?6䊮Ò����$�4wbb�0{�շ�d@��{�fm��xlk	���:ݨ]D���N�'T��qV涑S"D����f�H`�c{N��s�_��^ƽ�����&���Zb'J-�:PgY�������/�J}�L������o�����Qo�#v`ׇ��Ӭ��D���j��E��wC���M����0F?#H�����){���Z�z�A������j)��~#~��δ�M�/�A���Y��M���"�~8x�p��K8"5�f�l����2
�֌oj"�����,p�
ս��C=�*�k���Q+�F�O3�+�4�=v��P$�=Ic����Y'I �s�6�r��$=�(�ä��u�8dq 	\<�d�t��Ǫ�Ɋ-��\�2���~�����׊&�)�[��%K��BC5�&�'�����n.�Jk\
f�xqD=ؐH����o������A�����K'��H�ܬޚ%sc�����={��S��M�כ`}m�ΧqƸD#�{�{1a��g�yR0�U�:ßk��[߯ȋ?1 s�TT�Z��uL����ppؼ�_�Q��yݴ)��[����h�'�WZ<ƽktϭu���h,&�&6�d%�SW�UNf��g;ǋb'��ޗci�L���UNzϼ��v������AWH��'/Gu��$`xy֔�Su��'sMEl���+({0�����(�K���� �lw�?p�A�,���Ŋx���^�#�����)��;I�cVE�%0$��j��L[@����:�B��}�����j1�P�r�I
� ��}�����J��l�o -�\Y6a��}:��P0{��������3��wl�E�r�6���M���q?�Ⱦ�.@���!'�5Έ���i^���K��dɚ0���BBk����	��-�g�juY��iO ��ً��]G��9��J�Q.�]KY�<[�qZ�����,�Ŭ:����N�*YVx�1gOh���<O9�e^~�Д��x����\�v(���S�-�4���IIP��b�@ɏ��Z! �VU>��t ��_�>{��Y�ڄ�A�U��*�.g��(�u_{���Th��Aʹ�ݩs5J�v�+d�<�R���)��.�[;f1Oxu�<���Up��Uoc�E��޵�K�T��v�V���"���EDTd��|�٨��n��#z���^ߤ~ϵK�q�@��l[X�|H�mk�ΧW-	��`��4[525ʎ�7�Q*�sz]�J���������=�8��R�1j{�U�6R�fҸ���Vڃ�zoS����'pc��
�Ѳ�un�;����!��>d��g%`�}^	�L��2���j������0���3�t��Uұ��ҥ�|����t��2R�����z��|uQ����q
o���̢u��F��$�l\3�a7w�lJٙ]��=!4h�~?�f��+mC����s��&�C��-Zj"{�V}d�E9�+T�R�wz j��c�	UbX2%���%M�BJYA:�V���U���� 	�`Y'�!fG�)~����n�u D9W%x��
U���ހ��NS�����`�3�>q
b9��;�?"ԷVz�u$�YB��s{��67~�JJ�E�']���Ie�->�b����]|ч-�}~h�f^
?|��^���Q=JQ)L��;+�;Ř�b��+WX�Cg�j���;���-��/���ʉB�)��W�O�"�✀N�C��(1����M$�5s�bs�'`x��E���e19�������!�D5�����}瀞E�1�!^�S�{}��C�f�@d��>�
�(WB(;�_v�������n��=��D�9�3���3OF���7���S�eoib�Ű�2*'9��%.�we.\�A�����j_L�⾖��Z�n/%�����P{��;�A�)��pܣɆ:���=Ga��u��C7I.z��a(��E\�r�-�m�Cb��'JP�pC�'aB?�H�KH9�mv�l�k+ʥ�.b�����"�g�7�WZ�햪��"�z�"+�}�=�3YK�Hͣ�R�����#�^�T�Z3>M���N��ɪœ��Pb���+2G%����8b�Yc;xԧ��&��[���o���7�PW
Rh.��Y<B9�ǽ Y��#��5��s,`u�����p9D�Ď�-۳��ӑ�ڮJ#�r��!5p=0��31�a��ȿ��-����[!�P�s�V���3�L�ϖ3�"3��>.U��$)z��|�Ͽ����%k��Tf�n�,�'i]sU4��^�ۑ4Y�:aB0w"c�ْ��;E� �d@��qY/��W���G�i=B=NZO-��f�!xfԪ)7�'� R�U�E�Gm=�A~���\�2�N[�n#s��,~�6(��
�9�3�-)ѫ;2Ȓ���l�.=v6����>��!(l7[�b�yy6�/�ģ��}F����7�!'�]`��׎\Cnv��QpcoTsf�>9���ؿ���u�T��`s��D��`sʊ\�Q�tV�r�{R�ߨ,�t�W�zC�>ߝ�e����	f���m��A_�0C�&%5U�'Fj���SG������ȕ4�[gj��>ak�FX>Fpۋ�N�D49�6�����d?����'��k#(rO�����A[L���O5b������"��&WK�2�t�u)xCG�7� +=��؄�����*%�`�����H1B�	*2vO�o��Z�Al��!k��I��l�� g�;�1]&z���S9��;~&��g���D����ܯ�iQ.0=L����V���`F���QK�#E����B�Q�c�}#B��<��.^��|lK�aw��R�>USf�䋬�x��y����&�@��8m/��I���-�j�&���цhe�-�d�8Y��o�4Q%Sb��5m���o�h��(�pS�3!,Y���&1��꟯n� �������m�&|��Au��%�����x�� EJ�{we�.��-t�.i�
}4Q��`}=����P
9ފ�������^�����~�z��:뙈��@�2g���%r�t�ͮ� ��.$`EC�i� 3�6Vo�ݔ��"[�.\�d�׃���6{؉ 3�z>�#�9��w����V�c#6�ݑJF�s�=���E�b�g(\�(u��fZ�|���{Js?�ظ��/��`��]2BО,{WK�qd�NR��Y*sw=[Y�"�VC���g��3�M�!�^�e���($^ZU�:3C6��9W��n&�g0���t	h���7HZ�zQ���%�͒k=��J�f�h���\M��:QG�܆z��co^§��؂~#�̪���y�. ��]��o���8d��X��V�^�R=����y���,��qտ�<���ݢ�8�kd�������@"yu󋣁0�w����迳� Ozu��4>���l=�?�$��!��#եW���,�*�k:��+��r�G��M�`fή�W@�j�������{���E����[&N���Yq�����^j�v�}�Z�ᘑe�n�h�l��K%��9!�甁�%���B&y��Vy�k"`L|��9�`6���W��3.^8? �4�����̗i$x�*,,PC�2�5�J�d=��C$7��Fb��*��LB����j�H�_��N��NJsRq����鮡.���ya���+:���,�Π�sZ3���(���T�J � �R>��1?h%u#~TώfǢ8J52!o9���(�H�ӠNko$k�%v���Q�%�F�6ì+�̂�F���=�5�@�kbI��J��?�_����E���p4SUX�g���^s�$�0��'�E�7y�@�0�A)��O
�=���qoG����v&	�iY�� ��CK:!q�e�S47���@���dZ1��4�0K��`�&?�����N�#0��h���1�c����DS�
�4-@��ɛ�5Eh��Ӷ$�{�eK�z��͸i�w'6���M�E=��ku�l��&?B7�6h�Y��S�҆�oS�#h����UO?tN	i�<f�U�;�F*�h3B����I��f�9��r�2muR"8Fy���%�gr���� k��:P0���D�(�@�����S.�a�_��lS�͉�/ M=�z��,J�*Wei��τzcSY�o��|�lP�`�/O��uR�V���?pvU�S��D&��&��n�]oM��U��rۯ�4)��j;�r'���U�����\�4�txT��,~:! 8Ye���Ƕ���3>+�{��7ӥ��\��Wxᶚk�[zV�f�k����uc(�&��d�&scQ�-ܷ(t��L�k� ��
��U��2qd�֦�V�q��A&@�d�Ec��=��cE���Mfmx�vY��Le��dF3;:-�Z|�m��oں��y䐦G5�֘J��8�?\&Թ�Mƻ����a��Bp6G��z
�dqI�S���;�}MwPԞ���	����;�B��3�.�PSL>\V�5�wv����B)d@��X�!ͣ��`����T����]���,O�� i����3x�����3�B�A��;@�^��Ы�$$A�џ�T���pƽ2T�L
�.���]yr�a��I֞@	�i�,�^U׃G�+�L�I�ak�\`� l	�����