��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&��n?��1ů��> K�-� �&�T�Ek/ֆ�\�놭5�DꢘP���+L+X�4��J��#�0�8���������l��jT��+�(���������6�MC!D�;�m�퓊D@v_p��䙋ⲝ��C_�6�Ռ��#�� ���	RD�4D��畓7���vn�H���0���fX����4 �CS�C`{��;�L����li��� y+����FD�p"��]���y��R��K�({� .؜M�������	^5���ɋ��&���&�@*���
e�� �t+���
_6��O<��7f�M��u���m(MrN����z�jL���@T`��M3��c�uQ�Y���%�dD���,�~^���y@Ga��(����C����	��G�86�S$��ɳT�ز8���:r��/y�[ݦڍ#A�����i�&<nU��<[5)�Z�-Ĭv���0t���d���"_���:�'-��d��*��q����_d�y�N-��~";#��������Y��؆���	6ZJnԷW��έ$Y�K�?�4���L�w�Wmiɶ��Y�?jx#*�i���F�m�E����O6T>]i�_�9;�!(��kH7�OS��_��[-M�((��lO�s�$�g�x7`��ZV�E���F��,9�j	@���]}<�ahb5~ãdl&I^�	v����-�@�@���	��!��d��`j[Q��� r��;f�i�.�m+UH7��/OV��c��������l��i��M��*'��?���G� SK�M��H?�ç��q;��)��Rȩ�"@���r��Ml>8!�S��L��EgeH]�8��>]GR=&���C��i�Za�z�,�F��h�q��^���wT�a���%�9�n��?~SИſ~�mu�OlIv�4'sT���/a��^��9��*��G�Fh�DM�_��CN�<�_Pg��O5��}s�%��m�o߫R���X�Q?��dK�Z|:�=��yo*�Fn�e��$��"f�$g1�B��IQ[��M�u�?��t
#�&��1��[.$q�ݎH��� Pi��c�U�U�gTZ�����i.���:�����Q9C��?ae��lzn���W���5}�`:�)������$ہ��s���'i���q�Q�`�<� n���1�4�bF��9��f;��>��8A"Ʃ�R��0X�E�=Q����|�56�V�H�����-�\|ڡ���٩{�$�k�ɝ�?a���pi.�uE�_qU��KHm����e�u��Q4�#��
�������c�Q��XMv��2����3s��G;�mH��ȥZ�s�y��n���vqYAy$lM
g��{O����hڰ��c�u?B�=5�Q�Q�|CM[	�SV�`@`�o��R�Ȃ�uά���ј�O��Ք]|���!P(�"���/�ӈ�TP�	�h�=��N��8֦���F��"���GS;�F��FP��L�m�ʠ����Ĭd'�%����֨��Ԛ�� r/%-wdr�Ҁ�O7�v�"��/�� �4F�R�(:�ڱj��-I�Hn�݀�/J�[7ţ�0A=���d �O_����������+2
�z�I��pr�-\Q�JA��Fc;ؙާ �(�X]~?�2�&\��1�W� 4��F*Co7�]������2�oK0�=��)����č˘�O�t�q�5z����<I�D�ܴ�6F��Pop|��d˳b�<�j0~4�#&�Մi��ldz�N�k�&h$$ee�V�s�n=� ��#�R�P�r"���>��]��I�k;�ih|���'Ӊf�t+�45X�o��	��)L���TikhN+P�Ym�ČH����w�����ꢫ��H�ҍ�!��ԟO܃Kv�V���J9��@?�rj1�i�5*��#ӛ�}=��@��c�|�D&[~���Ծ�b� T�Iq.C��]���p_&JW֣w�d����f�R�_{�o�_mYw|���i�g�������y��l��S���n�d^il��nD��'��\.
_��\�}�9n�N�Ye�/&r2�::^[L]逷��P&xj�&t~4�P�Ѓ�����,/�\��.?�2���@������ ,�N#�[6<�-�7��*}�䑤^��k�+�0���5l�38\���uj��^�O##(���lG?���#�>�1�:RT���J9�By*!f���j�K��02.7t��l5Џ��}I�D��#˃����
e��p&�XH���67Q�.C7�y��j��=V	xV���_gʉ�h�cD
i�-6?�9�>��ϼ �����5�ݯn�loiL�����X�}b.f�z1�z�Н�����]"i\{�S�����̔޻Ew�'��+���3�$���I��j~Xc�3���Ӧ�Z��Y5�~p���"�+W�e�(��^�Ԑ^��^_��K|�Y����K2!�9�H�eҋ&Y�G��G���^��(�2��/��Y�G��Qϟe\�w��U\l/���9����pୱ���e�$�w�ŞK�S��l=�n� %�v�[�}fȘ4_<��ꁳ�M��3�)C�.3F��p�{� o/��K�����pr���"sP���e~"�<�1�s(�m�H��Z2Ur5j{o���e=�����%��X~�����)���s���_��t�G�����>�=�IO�>�
�ο��5|��2d�q��JnP��\�B����$�sh�ؒ��p�#q�7�}W������-�1>)c�f8���1�mX6�^H��!r��}=�3��n����m:�����(Б�bt��,q!c@|72��Q����pU톦����l��O���1���@ž��G+�q�t������J�6z?�A�c)8�nL�%dͯ�s�����ނ����5��$T/e~��'��"�y�^9���D,���j ����3�5H��۳$>�j�Z���M&l��yI^��@]�&��~[�Լ1`��9��
e�%��O{_�E@
��a��و���5�
�|�`	�i��.Ҙ~	�4XF�����e����؎t_���I��9a�	0��)�q�l�58ȧ�#�W*[���ɮ�Ü�?��/m����bvb�x�������i�N'o�ms+����v4#�jH�������b��y�xeO���,�X>�&3i�p+��0ŪI���c�=ݔ'�'o�?�bbg�5��Ã>&ȑ�7�o&�q�[6�R�����14 ���� ,�klE(��<[V�_�9C�����m�Y5�����ĵI��W��ͺ������>�7{V���d9E���.��ڢ6ۏ;�0�>��*twNO�D֮����y��J������Qp�����+�i��}�9����F�\Q��ʭ5Nʈ{�AF�����4�6��
���q�f�aG���>҃�}����d��̫����pg��ʆ��p�<�H�_4猊����D���3�����f�E�P��K�"gl>�)ד~= ��A��;�j
��8�����B�*D�a�ǰz&Q���Ti�eqi�}��B�0�_|_tCa=X��Ar���P���)g�E���~By��pGY|��a�M�� ÃX�b��Ѩ4U�o���ft�/� d��"䉈wY(�.Ŵ��4���ِ�o�*8L�!���Lz�a��n��b�g�����f�D��ͳ����1���_X�
�N�C��0Gc���U~m�nH��٪
j�R2	,�h8��	���*�vP<I�qCs/L���K�����-P<�(b^>k;N��n��^�҃��a���*VQ��p�?���@���F�SS7��"z6kU�mE���=ʘ��R���y4:���:&����xk�@j1"Մ�U:�3�V�����ߓl�$�� �oG`�p+QUM�=�wН�@M58�<K�e�W�%�	�Zy&�T������׌��3T�ͼ���<�Js��f�5�W��R�����L�\�8�Xm	�������rˊ�m���~y��������F�*�C���)�� I�ٶ�0;����ɛ�!G�8	\3�T��Kb3�lЉ�`��&�n�s����һ�F~��oڑ۝9��ۥ�9�G	9��Z>H@��Kg�*R��é�]Q��ۆ�0�2���2�ha��etYx�xH`�F֪9l�U�� ]O~c?��֓IJ�C�)��w�[�Yq&��n6����F��*=�L�e��R�f,Fq��/�����0��N�J!����am�G��<�2���_�F�V�̶Wz?`� ����Х֜D�� q��%�~,�9��l����	Ε}�g����0!N����fR��3�jT���$��P3E�T�ǋ���ь���� :��)k�;�z}o ��Y�0�;�_�������[嬆����/}V�!�ލ�/�С��#n^�	/p,�ҭ��`�_q�j�b��` ��Fۅޢ5�j`�e<��w�<6�QwK �Lž�(�����?�jLԋ[�=�G=A��A��˲4Gi�d=���~��* @��ᑯ�t@�ȟ�o�e�^O�j4��O�MA�	M�4@6�⧀��%�.����r�hқA+˘s
>����l�� r)7u��6��V���,���iL��A�ղ8$ҿ��+�9͛ӵ��3q~}ymX�'~����_�F*��?�T�~�]9���bQ�N��:�ti>��7ve��$����w#�i���3/�w����6'kW��G!�4������^������b��p(��P��b���ݯj�ç�
c�P�j�2WzX��N�<RОO�=PU��X��z����I��^@�U\F���h���x�{5PM�Upٜ��ꋥ�?��灕Ŷ	�C�?�F�.`΁���a�ҾU��,����<Ip� ��_��z�).
Us��2��p�Z����*F��Y��W��FH��E4�guğ�m���ꣲ��͒����J��]�]�~[�#C���c
QC���L�>�/vgY�3����ҫJ�3�|�Nd�?��/��vY,������ñU�n�ٽ ���ѩ�2����-O����;=��c f@*�>M8=k�� ���>�|yj���G}��P,�չ0�sʆw�R�����+,̛u\Y�����oz&X�%]�'f=�h�Fc��bJWM�4n4�Ⓓ�����y����ω�V����GV���~��3�����������H��d�J�P,O�W,��(��̈́�p����L�W[U�SK���s�E^B-�XHBr�5�a!�ԡ�P2g�!u�_cw���@d�`Մ,#e^W-��<d-�Ah����:�(�h�-���x��~u/FĖ��,u�\��\��?��)�6�A�^ʼ�<8�CJ�]�#f�r����
5AwTa��u�n;�@��"5rZ�S�DS8�kgF0���s��7�����Z�/<��FP���x���+�`��KA1�Е�蕹���J7��|j4!fU}H�����Ј�pB�+�Gp=η�ؙͫ������Ř�SH�u�9���MtjC�mߎ���1���r��:�����6�����\W2�g&󧡭�
%������v("��),�փ�?bT�x��� �������濴��t~/[�̾��&�ڰ|(���{��^���r�R��#@��M�	��}07�zcR�55��?�|��0�Ŕt�f@�BP
�N)4��}�"Al�����L,��A�'��XŲ`*đ�"�_�Ff��p��:���M�����^2_�Cp?7������#鍑���X�eb-�����j��F�ӟ2�����z/O�RE��,*y� )�XUt �������x�fK����d�dv��]=C�$-�	�g����B�wACVEj��#��Zxɭ��V|Ꮵ�ON��>�z�23o&��N�x���
�@�Q#��k�{���+�>��X�P���]M,���j� �>#w$�6��bpK8���2�ьJ=iY�t����}��.�t�;��1��垍��	W"�+!�P��.���8NG�<?����&ٱ�=�zl����n���p�݈�b3拙]]+����6��SD勫�1�t�/Q�ĝz���������>�������Ǧ$�_Wa���9�(�U!V��>J?��,8�A|�𯫑�ǔ�FN%���yK�֓�W��bv��ƼԽ@�>��-�����b�,��q?�HC�R�S�)=�^��7�ȅ��򯱘��N�iOU.DaM�$��$�	�fر�">�>.N$�3|�7�<q|#P��C���{O�˔�i%$�2�Ev��|ܵ��������-o���OdǸFv���XQ��<0to�>$5�ҿI��8�&�W3:s'R*�|[e+:��f|{{�.`����PH�1��p�ov��Mx �y�&��,ea�!f����y��n�@R aJڭ�=�s�.�E�}�a8u~�A.�爭��5q�S,ˠi27��w�r�O�|���(��p��:�r0������@}�=�������-�:�ntJI�#��}�c
W��*S����9fd0��5�PC��E@�`*Oԥ�sy��ȳ=a`0�t��4�0�m�����%�9�@TRH�b�4A�8����
al�U�i�����u�oT�K"��If|D�s��~�Ic]�9���u�uUc�7�MWP��K^|��,������Q�)l�O�\��8|���sI�<�$Tx{co#+_��I/�n�N?t�o�@��L&�i�(�^?`2�E�L���5�<O|��,D��ɈU%
��U�<x�.1<�����ȕ���[N5�e�yC�|Jr�K�uƑ1}gx���ǎ2 V��0��������Q%(=0������]�!���zc9p�p��[1�[{���N��z.Y2��fF���H�N�%��n�� |���������ę�m�8�-�ީV�4�^�`�a��N|��N�T���r$nL�]gP�.��˺H�Y�jP��>.�R�\P�:�F9p�Z�oF����3����&60�d��p��[��B�������lj�&ҫ@�R�Q��w�͸][�fkOEU]U8�E�\��j�~s�OJ��grX��+{�������Q�ȁj@� 6s�"��?jث�r��SԠ�<}�.��cx��(��7�)|cb�F2T�I~�J
�C�)E�BX�o�9��D�pG�ڌuJ����N���d���|v}�Yui�̗)q`�P�=�L���O�1�zq�a���H;���9l��h��r����)j��q�)�J�wk���PhPȩ�����$}MIb/V����j�>a3�j|�[�/ b��k �S�u�!1�6���ri��)&˂c�*�PB�"������Ӗ�.K��^Ȝu(�5�#*��=> ��X�SBw��z�S�W8|~�J�[�.'0�f'��H�;*a���J�(���s�μ|�o��^��x�H�0d��]���v��WSg�Aeg'fn\q�p^ph���TO<ZR�����$Y\w/f����;hE��T��x�	e:Si�W\�TE��E	E\�dy�}���%k �� B��!�ү�v����9�{���K0�O
�GWP���ŋ	���+��Ǧ�̒No����ŰG>��V���g�NcsW�2�X�u1��w!:磮E�{��l�=���#����7���<PhULrq4^�MԔ_d�����aƛ�~](������#����3>
��H���K��l�1D,FБ ��Oe@��@��7�x����yD�����C�Z��W������V�d�Y�0âfQ�-�] �1��FA�
����h���ֺ�� ���K�?,��ZS""'ޠ
��3�� �N��CI�}u�d柌'`�|�GJ�޹��T�] �;w�ݣyx���o���@M0l���zY���~m|-@6)9j)�?�b�g����S�"���<�p�E��B\���*�&����0��M�O=�#�Y�-�U&}:� 0Y'tAN�µ�����U�&�6��p�N%�}2.U�z���
�F>^_�<�S����~'%ɟ����KIP��M�(Ԧߜ������<Ks�5���D[�n�w ��-��n���z�o�+M�0�e��!$�x=�N�޶%Q�4��8rup�Q#=P+�~�*�*����+��>���C/�(�c�X�ɑY�����R����q�t���l�ui�e��(10ӯ���T���8��	2�B�9|���꛿�D�P���݉}L���n�	�B33n�m�c�+߽����
2'��*�=N�=JoH��(eX-^J�|�S��PZMs`[d��	Lؚ�W�!�*. q>����]Wn�dG�~����뽐g�L�Sr|=�IJUM����4�w�Y1��@�~�S�v�j�����S�D�L���g���Je(Ǉ��x�J�/�%'EŊ��%��wX@���ʅH�'),����)��H���T�P�lƺ8�PL�����dN�o��>�|���ƕI�h���!Ҙ�=��������4�Ȣ'��ك����@(؀�qYig����;����ʃ�O��}�ڑ���FE�{�r���G��^�!4"M�U�	hw`9Ri�m�E�s`"�]Q��c|���
$��1?L.�����809���|ֈ}X�����N�l�n�(\�����t�SF��`?Ln^�@0ٰ�ކ٢s�O�f���{����\�v���M�ٚT6����b/,)�|�d���<g�P�D�`	8�j5�0��n|�+�0o�-���V?�&���G!�8��l�R�G�=;�a�|�ͥGP
h��3�C0�m���A�����<��ݑ��YčU�~"���K�x��av��{�5L�����W���.��HF7Pfe��CA�#�g�?�Ye�t��yġ��GsXha�n(c.O�.�����lN-x6�G߿i�r��ԍ�L�J����^Z��ģϥ�i�N�P�MYB�͓S��竅o�Q����-�����8��Y&���f��+��sҿYL�^n�h�q��:��0R�l�R������v�&#����gZGS�J��\�B���[�oU�F�_R��䭙�����f@_O��>q/�8�������^,�e��_468�M�P8�(��53���mP��Ӏ͘�F�P�Z�%�Zi0~�iF��v]��ȀCt3�lW��5Q;Z�bl�5�n+�*�������[���Hշ��Pr�t/�ų��?�����u,X��K��i�uj�L�H���L�F�rr�܊�3�]�Ҕ�&�'���pp�.L��~� ����u�̚p�} a7��C����P��{H��cv�8=����k���:me��k\[����1�}�$Y�k�5��|�!��9�z������+a9j����3B��'�WK��w��{��oB�b�˗��+��Zc�r��7LLi W=�\�����x���%TC#�����[�SE�O`.�Y��XCs,!��[�8�h��a�/�u�����c��QC��_n��K��Ԃ9�|����I��i�bԃ�4��O1DCF��3a�vN�_tf��p�p@O�!��4|!5�:�H���<��>F�[����,m���qc'ڟ7� ����AO��D&?
��������#�a�oYPƱ�T�NcQ�@����O��U(�@i�G]����gU;�B&�S�-�dXa;n5؃n=��u��!B������1�7��Z��B�!���`Ɔ"~�osO}��_���8��
ߤ]E��b�+[Y�.���ryp�x������7p��L؇�ph��y�BJ��C��"��X}`�n�n�=[�}�yB�hu8o�VEa	�"XBPk۰�QG*�yrk�k�Ad2^�oL�� +����HP[�\b��m���H�7i�F��X�f\��G<dҁ�K��h��s�ƬT�"��.�L��p��#ֽҫ�I�R9"�/���t��W��_���r_����	\�f�&ICP/��
�'�ͻ��cZ�Y.c���kɆɍZ�I	)Yl��n�� ���d��� Ne���UY$"��.�)��a� QR�=�\?.�j
��P�)8��]���f}��ڌ����x�.�����;��ce����3�ܕ+u���Gv��#p���ȹ������W��Fl�V$�<τw��m.� ,� ��r0廨eZ}P��A��;��h��y��7*mBCf�n����`�t��h}*nfkD�,0/u��6;,���\9�_A:�c%Q:�TKL������g�M�p�{T{��]7��t XQ.���:�W�P̐��`cv�U/-äCV;��
��b��e"��)����i�It%昫ո|c(��� �v@�S�Y��ҽk��z�f�3m�ٻ��ǈ�q�ԑ`0sSU5kv0r�GW��e�����O�do�"p�o&�xj��^M�~j2�C��Cu�齫q$��R����*�W�_�����"H]:D&|l")c��+۝���*��T�ţ*j��51ѩ5�2�!�*z�Ү{9�\�)��'"7@�@+���Bm�%����H�5�a�X��������߭��N0dWڪ�ț��f�SR������WԲ
�/~��'�i/�F���_�{�B~>�~����N�¦��gq}�v �<��
G`(r��8iR�G������d>���(��vnĘ�:�߈SkgY#�$�D��U_6	�D<2���b��2���;�
$U��zmu�S�,N���J�,7D�qC���=JI�AB�Q�y����
c�y}`�51u�B��g�~�Y~j��(5,��y4�(��+p9��e����_�"����z�V�!��kJ7$Ɗ���Ƈw�H�(�n��G��1�P��ug�g�R�+`�ڭnP�9�0*�w9R���Ddg�8�hqnެ8���* ��O)w$���SBk��N�H:di@�����y6������`�J�}��m�F����+\����=��/�h*E���#�<���י������!��WdR���	49�T;�g�B���m��5�hD��J	�q��"��&��yA@B.[3l�(/��-��}�-��5�0ѥ��W"����(�a�kq��b��N(ΙA�g+A��?�*JEm�����N�l��R}M��e�*��=TiO�. ��U\5V�	gy�����~�^�ӞW"��w�U���t)XDZ���\���&��yƐUn�c��b�`V#�6z�Hjy:�U�/�8�A�"~�-G�����Ǩ7���������'W��}�*�Xk�-J���M�ӇE���O��gO�
LgQ�$�fT����a�v	>�
w��v5bI��W-}6�dK��Y<)���"4�DY��n�f������B�u��^��MըE905:��Ӻ4��٩�(�}����jL�=�����wi6���!z��</�x����bTچ��oɧ�.�=@C���iȶ��c8���?���Դ�N%#OC�Ȉ�O^�L0��6���e�u~$�YY<�c� ^07<D��ȻN`uM+������0}�7������g���)$��z6���-s��P L��Vz1VQgb�ׄ("C֊�@=�h�%<������@JZ�c�[�M�`;yf�:��P(n�Wu!֦���SѳM���T�g�l`� .���٠t������]�;o�Z��~�ZS�g�P�n��q
Ywc[�� �c[���N7��׷Я��fp�'?�x��-GQ`^�D�pK�����$��gש�P��k��� FN)�˖Y����Ǔ�0봦u� ���ݟ�7�~2x\����"���)~�^3�/t'�&G~T ���@�t�m�wl?������p�;!OƤ���پt�d'rYR�-��!a�?��L�3�\Ө1ah��:����u�P�jMQ�,�ig���˖D�t���=+'�J��T�y��Ғ�ŔE6����e����]�S�ș�8�rg�T�U�Y�-����#�.����3ds�h�����R��a��iԓmQFh$�_L���;�0���y�`v+$�o���*����n��ܷ3~�15dgt�?�È�x�����(����P0���k4�v���B��'D�CeL���p>#��= �?K��q䬌BÆv�
!�u�����җp�n~8꼃��L��1�3�%M���ĥ�{��'	:Ո��d��g$<e�2	PYi�(�k�p��5Ք�ۦB{�'AtVo��G��e��-�X�zXC�`�q���SH�7p������PI X3��o�b�mm�VE�&�PW�.��:�� < �XS%l|�Jܣ�IT����Z�{D��,}b8k��4ft���3!�ز��eCg�g���Nv���ڪ�|8�hǝ]6r������/O^�f 0��g����P�W�uzP��t�c�\�K���3�:��Q�~�V�A;���m�l��U��U���"��J��� 7O�E��G-��@;����BKo���(��.���k�ţ��L/@�@��F�x
m��q�\���ZS ;hXj��?LLzgsc=�Qc�j������/܋�ke�g����lN^&؇�-)��n�)~��w�6t��*�S96�=��rQL� oϛFz�D��c�a�&4d����83���#�2 ܔ��$���Ŏ���̀�{�g��9K������.̏�Qze/��C�?�̎�{"�A��ITz���|RQ�����.��N���5 ��7�f �k���B�Cu~�n+�h���k�b�T\@���&�Á�pp�{�$���y��^�0ς?�.ZҮ-
��L�6���z'��-;j��L���]IC(C���c�y�LyP���ly�CH�9�o1��fb��Vk��y��Ҡ��"��5��1]��0h���`a��HR��ݳ�g�A7���fǘn�$�1�&9\t{��钽a%���!��b7�x����/�┦eXv��$Z�]nq�&�E�F�*o�5!k�0�������Ѽ��� bg<?�l�e=�\U��|���@�Tt��c7����E�,��3�����!�2$�!��nb*/ 5���I�H�*O�:����ɂ
Q[Q��Ur^��~4{���YM_?$b���7[�0M��6�W$s�NN�O�6��"˃�u�	�D���@������bA��ZӋ+�����V(���TŵKF=[Ã)j��#�	K{�P�u��e�J۝���� �Ď�g�NI�y��������5��gK��Nn)C���f������ĚF�f��[�B;0��2�(�"_��SH	`�㫵w�fm�/�	���S�(�}-q��D3��gy�e?ZlV�vyh[���:TOo�A�n�=PX��LB�V�݀�X���[7ԧ<u���q~G޳dC*6��Q[�Wi�PG��>:'\�T#u��P}ұ�1�<�U|���TO�:�_GV��_�Le��5Ř�ռW!�E3�'���vw,bڙ�	�d�E������[p�ܨԝ���sy��o|����,�R�R�KC��L� ")�<��p�!����Zuz��j���qp���oWb��?:�>Z!X������3ke\��R����6���unl���v�׿y%C��_��eI����V7b�S��=�pj1��m�+3��������i�3]T(T�@�7ץ�0���L���\3�Z�o�<Qv&#��K ���[����X���0�f�A�߾����Ǉ�g�����e�d�FX���E!hr���H�M8���ql��9��N[,R����_=~F]uU	���@c����E(�����BTOB
h�3W�^�Fl���c�X���	�1+W�M���(��C'%<8�O�ٓ댇�h�zH1�E����[_S��P0P�{��?4�o�`O�u/-[DG<���5u:�C�oS��b��YR<W��e�(�=]�#`��*d>h�q�!Z3ka��Jc9{K4#n�AӑՑ�Ł�*"������X`�����p�2�}��-60���������\�C��x߿xU���I�wͰw��^hp"��L�y��sK�J��OfX����+�q����3�A~�T=E�'l7���j�,�*#b�>�r�o�M(VL�T��v�Qt�-榄1�?��8\�Zo��_3�o]�~�ro��8�M�����W,`�$D$Pq|��I�Kb�� ��D�\w����>�!H1��<}�]w)���!<|G���3_��Uk'��wp�/�L�-��YgM������{� ����U�s���L7��i��AxK�/�F1�[�����ȍ��ת���B�����֕�+�.gX�!��8��Y�����!��ݵ�%�f�J؆���1�Ј������++�ɱ�b��J3�B�W�wm���J
�k�JCT�j���R���FP#��E���b ��,�����U�	t'w��^	����b�8)�����[�`�������d���Kq�P�ӗ������e����4����D,�}���L�2�{۟V��9�d����W�er?������ŚVq�_y�5�z��/D��ߟ���ʒ��f��Q���,i�3�\]�N��]�kۈ��*�p��t�^Ʋ9E��wL��8ڛ������׋���3{�xŗ|g���V �Q��f]%�c�+��ň�"ê�4��?�5Ô�7.�s�lH���[_ߺ�+�߂���R�e�(L�I	`��E^r=��+p��ܩ�P�+3i�$�����08�<��XD%�P����9�gyS*JX)���Y�xi(O4��a��e��eL�ѓ*��"$n��t�(N��]I9��Z�i}�jG���?�K:��+�<@�&�=m�-kF�7�$���^�Ԑ�VXU��lT�G��aL����U����3��w��3��_���qnP���t�R&g]rE�rKh>�'���ih�::<�j�마rB�4yY<}6���G3pFY):�;�҂��+)�^Z���J��6�\P�"�Ⱦ����a��[�=���b��-�Ow��|��Aiuan+ݴkJ��`��DhT���~jeJO��� ���z��"�3�}�}�B�êku�S7���%ȍi�k89W�)��Z�|u���5�[y���;
j�����Cl�#̘H��=�^�k+|d�^�2��4�c���p��\2�e��I����lR���NܷY����^�Ĉ�����u�%Tư�9_ڪ��)���В��?rQ�ST)3V)�����r�2�,`D�=�p�ٵBV�<��I��55�׸�B����{�#ͻ������,CߗoBZG�ST�[��*�Uuٙ~�pX"��[(��$�)t�H��\i�|6�"��s���m��9�
y�Rˑdi)�'�X��	+�����utR2�~Ǐ�
�m[!a�{�`oPpm�� *�qL��%�`'�~��]����֥�Zl�I��#rI��)��S���RaIh��Fer���O9�|2��}ངJqe[oP�0|;m��j�s���[M��I� pM�\��M7��g�kٸ�B1}�|�pu�#�z=����l�M3{��G�h��:@��hH��=Dw��3�S�&�w�8^�3Tw���������&��{#-���i@Mj�
��ʍ�Y�|g*v�M9L1���)A��.�:�Q����L����B"Ve�K��Cx���׶�-�����i�� wxt�֒�n=]]ބ��o�Ɇ�>��M���Q\aӝ �&y�w�{���B�3�K��}��;���,�7)�|�_so�'���];:P2V?��S�N��c<t���0��b�7㵑����1`�`��i�'"m�ܧ��Lu��͠J*��p[	�K��,,���M��������m�2I����|'6��ǀ��~r_�~��
�)��$�( ����XA^~�v��}�:��RA��&Y)=��Ih �*����ΜE)��{ê��r�v��w��(F�L��Ô'�5�*̭ނ�1��(���а�g�P�����FK�f���mŀ QBL���*󬢖ɍ�����^ڣ�Ͳ�Ҿ;eEK�]{�sjop�eu�x"�"Aj ��C���xj:�t�(仡C7H�e��e�z`_|�@h����d-���v�<�4�-�:P�rDߩ �7S��-y�y���gB�W#���w�.X����p~�c����ڔ�Ƹ��}���
aȭｲ���3����-v'�
嬏�~�|Y�H���Wl���Ϧ�j�a�]��w`hO�8��H������X���N�
�n>����aV���X�\J�ه�S����P�<���t�.e�F�ƲWX�C�Z$?�, ��d)�R�K�D1�
��(��]S��:��/���%�j�^<o;���e��PMm`�>(Y]�ӯ^W�oIFY�n
.0���.��î�]�U1�����q�hx���,"_V(<eJ�:�q@�bףO����z�/�)��9�Y[���<K�d�[���a�z�x�^U�D�O` 6�*���A�����N���9�~<��l;,�k�5扐�<�~��8��`�C�`� ]	��:@W��(j�e�ʗ�28��Ko�ڊ��B�
��آ����I��Z�T�6D�3Z��#S���.xȴq�2]��L���Q�=Ǡ��^Fڒ n.�2�SLOx�{�U��k`�#����1�M�~��"lJnj��i��\��hˤX@��"��l��ɘ��Y43zA�«*�����?��]Q��5 ��^^C�GVAv��!. $��0%�m����?�h
�TW�'��d�?)�B1�.���y8��\���A��}dk���iq��H��X�Jo���^>���~})�(Zt(e�3Nދ(2��B�#mI�c� +��G�f
x��3 ���l�8�P��P(�B��B'����3����>�^��,��Cs��:$����S`�������u sa#�������Ѝ��-ٶMvR���m��	��q�%8??ߍ��x���E�a�o�@������0*��h�7ε �9M�B��q�c�iY����n����Y��]��9�d�r1���t.I��ؠ�۾7v�?���1�׍
����Û����n��B�(=�kۿ޳�[͚~Qg|L�jV�:g
4���I��N����e��.Sy~��kIl�p��"�����w��*��^��|����_Ԁ��M_���Nʘ4gnv�U��/����OJ�R�j=s@�Q�)MI��O��t��[t������ ��̴���v�Q���+�!�!���׵|��
p�)%�M4�¼��a����秼9�:Q/��m(K=f���c$D[��!�b���oK�pn�u'%h�*�<	CHq��xر��BI#��Qm7�<�������)�U�h�^~h>�:�'��[t�ɅEP��^�k��L�A�(Ī��|Cߤd���G��%�K�e;�Ji�ფ�j������t����Br�mY�B�&Aj�VHe]�6{��Q/6�_U��?6ܺo��a�UF����G�p|S�F�.��a���9�fe�0w�����*�ʤ8�k�`8<�@:Ш���Z�S5@�*���.�<%�����u|]+Ue^� ����/�R��|�IŢz���_��|�F���L���u�F0��a�OG_�����z�W�`!#��mUKqoHa�O�(�:y��CR��+H�^�6.o���-M�|���a��\��ݘ�8�Ws��rؾ��v�:7�Y���V����^%�9��A�P��r{�qQ�SL�6�|l���7W�eуKa����k�c-�ZBU/��(�������S�͔�i6�G7�Z��
��R�.�An�t�dc�Püԫ�Fḱ���'�U�c����n#��[
+{�x����)T��u�� �[1>ڤ|+@�9W����:[����{)�4d͉����]�