��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&��n?��1ů��> K�-� �&�T�Ek/ֆ�\�놭5�DꢘP���+L+X�4��J��#�0�8���������l��jT��+�(���������6�MC!D�;�m�퓊D@v_p��䙋ⲝ��C_�6�Ռ��#�� ���	RD�4D��畓7���vn�H���0���fX����4 �CS�C`{��;�L����li��� y+����FD�p"��]���y��R��K�({� .؜M�������	^5���ɋ��&���&�@*���
e�� �t+���
_6��O<��7f�M��u���m(MrN����z�jL���@T`��M3��c�uQ�Y���%�dD���,�~^���y@Ga��(����C����	��G�86�S$��ɳT�ز8���:r��/y�[ݦڍ#A�����i�&<nU��<[5)�Z�-Ĭv���0t���d���"_���:�'-��d��*��q����_d�y�N-��~";#��������Y��؆���	6ZJnԷW��έ$Y�K�?�4���L�w�Wmiɶ��Y�?jx#*�i���F�m�E����O6T>]i�_�9;�!(��kH7�OS��_��[-M�((��lO�s�$�g�x7`��ZV�E���F��,9�j	@���]}<�ahb5~ãdl&I^�	v����-�@�@���	��!��d��`j[Q��� r��;f�i�.�m+UH7��/OV��c��������l��i��M��*'��?���G� SK�M��H?�ç��q;��)��Rȩ�"@���r��Ml>8!�S��L��EgeH]�8��>]GR=&���C��i�Za�z�,�F��h�q��^���wT�a���%�9�n��?~SИſ~�mu�OlIv�4'sT���/a��^��9��*��G�Fh�DM�_��CN�<�_Pg��O5��}s�%��m�o߫R���X�Q?��dK�Z|:�=��y����&���o� �бy+�|�������:��������w���97Pnb���?~Z�wB2��بlK��Vʽ��ײ�S�F`���7��C ���q�J<�+P�p�^�s���(�JĈvJ�/�*��ҪD�5��V���L������p@�;�,e��KC�����-�h;�Z��
~׍ݒ�9r�l:�dX[1��qDJ���rsy���nԛl!���3���u[n ���#%���a�_�t2��B��n�ֽ_�}i0��tvp��Ȉ+�5�,���4���. ���}E[�\jRǴQ��Pc�1�n�	�H���hE½c�d���&�Qfqp���;���L�`ɣ^���$�)a��k���
�fl�Q��`Rё�c�^B 63�٤�_������K���Ɩ��Y!�	<o�h�C��j1.C�5mM��(�B�!�UG��z�����km�w��f�b�X��D�$6|aךK�|Fm�񢝷Ξ���^P��F�{U}�9bnH��0�E�na_�J5;�5�+��{-���^���i�м�?��O�Ơ?�7�~��H֒I�}M�'��ѣ��[�ʜZ�>����=�]�q����rk�wwb�K�YW�iQ����'�D�y����2�و�K���>��Ƭ���F��`n;*�3 ��ҙ�M��]����|��)�:q'�~��Oө�9�)��Mae���\S�����tW>�9���R�`���Zuk�FO7\���cq��J]UP�j��
��%z�E�qF�{�˚�j��
�z��l|�p����3�����W�Kq�S��}���P��5�&����;W^�..�=l̻�Gm�LE	��̪͞M�����0r�܆�}PP��Gxc�CF�|f��ќ�r���;�{[%��A��Sb5��fo�:^7	sb��U�M���F�Nz���!x݂;�8�>���ȇ����!�d�M���I�)g���N�����3f|L�� ���0Y�}K����<�"B]���c,7,�6: �PQ��^�n;H�2�`���3S1��|:��%��D8�ơW�^�fu���ͤ�w��Gl��51��?B囻�N���ĵ��ޞ1�]���󡦻�ѝw�6��-�{HU�-w����+$x~��keUK������5_��-{y����ѳ9�]��+�!&�1���M�K'1���F���j��8�L�U>�H=8�ˤ���x��&��qAF�%P� ^*^��K|���`ÆL�>�w�\{�sϦe�ו Z�]4��Y�J�'|�+��+nt/�է��A'Vj|����X�`� �.�Ӗ8	�r��d��o2�#G�.y�ܨ�W	v���Hܨ�x�g^�_�O��9}��R<A���ˌ�^���"�o<��dk�O��7�$ш���=�{T�t�A��Gpo�F�ߗ:ȵ�d5�h����og?��)Woh�e��f�8|��h�����t��l�����yTF&�<�ⳝ��i�����=r4�>|�@���s(
��*\����R���e�yǗP�n��S�YP�9��u�_���@�{��9�b�C��������Ѩ��u�����a����NQ�G�h��J����CsR��Z�.�b�0��0[�[w,��3t��Y�z���ٹ0�m�Hx������#fNPbХw�;۪���qϽ�&��G��[���㕍/�
����ʤ��h��ڷ�K�vx;�i�4~���[9ޚ�KeT�K.�?³�"r�o����LӇo�,��U�����"�v���j^X5�?�m��`�����X��L0H�O
:��m������O��F����sbJ��0��G��r��[���zy�.�cI��M�]�~�
r+Xa�U�t[�#�|JB����V1���,j	S��W�o�yZ{��Ba5QO��:�f܈��e���ߴ?��{TRl]�����B��(_$��9�R��-#�����%~�Ε���@tQì/c��[v���!��u�SWiY��Y��a�k��c<m��G��J8�قH����t@tP��&�\���`?]��.T.�����E�5�Lp��q��k!0�TZ���h�)�u����=T#�q���߬�Z����ׅ�FA��.�d�����_f]��" �h9+�r��uì>�/$�!Q�+J�7�Bȕ���W���៸.|���I�4%�L�Y�R�&ltg�� ��_@y�뼙��]�6�	�a��:����֍�M�|*���ט���_����3Qsi,�x��T�t�IkL����_�5u�T�s\��]C�^mGO��5H�JE6���K�ҵO�"�p1���u�Z"���gv�-��A�	�c[?�$&Ze2BK��N�/7l�̀C?��o���9I�$`����i�B
D�J(�kp<4=j㓶R���� `���1w�h�DыU\�)�v�.�N9 ���<���^�����N�͌~lה��J��2��i��ȭ�X�)ۅ��w�箌����8�L�z��K�h���z��-�og>��ڟ+օV$|9>a#z$�M���i�d���YQ$�v
=��>���ЗJǹ����X%g�3��c� ���~ �]�`�9�+)d�����&��^TL��:̆"�ʖ�H�|P�k'NcC*�7�;���ı̍st��7��`��XQS�4���7����.�$^z�����Z����v/)kR�栂��u�s�w���lL/0ge|p��g?�@�E	�@�ީ����c;���J���4�]�_sf���(��]�`���V�����n�4)Y����+�~fJ	�2���%]�_-
�֩'}0=d(X�u���{��;nq�g�vc�V��:@׍����N2��u�n����o}c��\���
o�(��]7$���#��g�x�+,}�{O� U�g�5>��1�}(BG�� c��߾�SC�Q�Yi�\=)�9����w�z�f"ӓi��k�D�G�>�Z��\e�Jk�>�m0J#:� ̳�
+�QZ�u>��M���Դ(�I�}rn��{,���lL�]W�_��z��<������Si��ɶ���hZ�D&ǐaB����G�ڊ�n­g.�������Ð�.q�M�3�F�ގ��+�bi���1�W1�G2���\pN!y�A����#i�~JOQ���]�N�����]w4vp��+,��0�F}n@��cG�z�iH�����v,8�\��K3ĢOOHf�Yk{(m��4Fi^��p �T�~��섣6kѴ�&ؔ�A�a(�� M��i9��/�?�ˊ-�r&�j$��0�5�֘�h��!��~C����)�ɿ��sd��v��P����I��-s��鹾�@�C�]��iv5[�y�f��=K`�~�5��[w�)�w��ٳ ���f:����}͎�x[��2=>��v
�_p��p����ݺ�V���W�{ՙ���7�@
(�1�T��i��)��EM KW�fCMe)΂�D���ͤ���G��Ɔ���sbp������_ž-V4�^~
MI��2Ԁo�;�O����L >F,���ʔaԃ�4��M��۹)(@6r��;��D@Y{��+t���Wß��>�߮�*�%v,%�[�Ca&7�:�sx1�!�щ����
S��/4-��س���&���e]~���4�.ϒ4��Ɨ�-�ȟZd3;��پ1��N%&lNn��}���N�C%�\��O�ݞ2���ࣛ��KZ��0mf���d%�΅w�!��(��/@�d�	.n���R-ͻ;Q��w�����$P+�l��+������n)��I��C��w���z,nT�A�ٗ�����ͥ�n'�J�vK�<����B�aZ�
l1k)g(�t< �G�����l	p��b��G�CB��=tT%F|ˮ�^�\o!j"�� �a�J���ɱ��ܪ��� s4��y����WQ�v�t���e
 ?��+�ץJ��ܐ� &��θ�-��2B/���P�z�	�������=m�iѭ����s��T�uޑ�Ơ3��1)��}����[+ԅ����'l\��z��@;�qHٖ,	Ƒ<�{. �^�j+�f\�cM�%p��}��&�r/��L۳��Ia�����{M��";j�� ߠ֩;<*���H�_Y�gx����06ԅ3�Sڡg���HOy�R���]=���JE	2���%��9�#ȯ�[e��9������M��9Z�P��=�K�"�W\�ï����:�9���D��I��qK�O4�R7�W���l�m©w9���8?Z~����_�����ؗ�	J�G�"{W0�x�m>���ڤ5n��T
�1�	��*Ys�,ҏ
�Y~p�G�9�S�8�e��`Y8,7u��G��&�63���ݍ��:Ch-.!8je$N�(/Y��`�y�Q`)���B$�d]��^�������� ^.��c�z��[۾�"����Dant�X�+�Y�C�^tR�=w2��cޡT�] >Y�:YxȠ-	͌R��vt��SB�����b��C��r�������kJ��~�&e~:�����8,��"�	Fg��V�����y��V٥yU�"��Ô������o���Nט��,Sg��ˏ��*<��	b;���D��S�G��3��(��mM�wǓӿ�(C������7�� �'�w{'��
]��tv��8�6:Q����>��Hy@ZY��́���v}��Gbx����Ÿۉ7M���BHz�E�� H����fr�c�n�;�-�{�uZ���E(b��-�3��)�(\],��� jS`��lD���̻/vr��U�+4`�i����/�f~���ӊ�\xu��fW)��!vXL
p���� �?����=h�Jw�`�v�b(O�2]}�'��xb{���lQ��s�(��R��^'����r8�T����?6Ӊ�����V�aoh�%����H�����/1�*�7č��ʋO���IL-���R?��]��4�)��:m�����;v�7K�y���J.��%��
�L�O|
���VW�#�9�J�r"���=,0����m��cHQn��|	�Խ<�߁&HO~�7л.peD�/`j�S�r�ĆL�x�ј9u�����\U�RS��Y�	�4?�#�B�z��R���b� Gd|�������bPC���&l���6�7�w'����eޥ/���x@ �M�yv��VC�8�-�$!\3��1�U���U<�k>�Y7`�PT���"��.7��*�prڢ�D x�v�i��{�(��mM9RL<
^k�@�X���S.d�X��|���d8[Qi��Lj쎚,�f�_��3L~8�ӯ�[4�-��� �n1�*pKr�!@�����,���ZX�.a�Ww�����b�ؿ�,4�W�{�Q�J;�q[�3��3�Uw`H��(�a?DeE��]��h�=�xHG�4Ls~�6��2p�}4όm͍ZI@4{�kH�#K,������c��b/�_R�(x�_��Z+��������䓜3r�4 p^q��E��ť�.=��3^��y$E>m[g�Ne�u��sZ��	՞���Y:�i��2��Y����X
l�Զt����D�#�T-���M���2�z���ڪ���|�Ч�P8=�xMV'�/��,{��8R.}	��O��Y���e����R�w����9�m�_�����I8�r6&a�4�����:]������d�ei�-l��^�H��u|�ke�7?;��oZC�,���"'�#Z+��t���՟长ݬ��v��OXR� mG�h�n
�NoN�� ��/H���U����Q�]ѱd:̹?�80dc���[h��5����xQ�A+V��l��<����~��zj������[/2�	0�"'�|�78�Jĉ�s�k�+4����{�2���7�d�Fu�Ι�'ip���O�8�B�-�å���V�϶ ��?���ݴV�ONj'����?i�N: 7��x��'Kz|��2�0�����C-4q��F_*�?ӥa���ܘb��
���sO����Ӟ�/��a�۫U̝;k���U���ސ���~�	vM&�.���K�2�E����25+K��71!V.=��
���4�Jf-!q?�P�V�q�E	��N%&��ל݉�ϭ�6	|
y��/і���@r���l��Bz�Hm�e��(-��B|��7���K�tz��]n6�d�C�s.�'���s�Vۑ�*ʋ|xM8�,Y4�R8܁���ͱ1&��ūO�'�l��*ZM�'�c��:�:1{��ã�j��'��I���������	��yË�zY'Q*ZG�^b	*��P0�dYW�e����� 	p;�i=����=H�X���dº&O�.���\3��,�-7�]<ly:nQT_����}2eᦻ[y1�Q��ݩK�y��%��gV�cs+��@�i	ܒ<�Dl�[�r���яޮ }ݽom�P$��cЂJɄ1H��r��{���b�v9�x&�ѝ�kF��d�.ˀN]!�8���3ėd��ˠ�eAfg�&��L�Ƒ��6��R��������9Ѐȷ��ʁ�!�#�B��WWW�7J��^w�
CУ�a�ri攽!��o嵼��k����;���(��K��f�hf\��
���R/L J/���UF	a�qa�M$ͼ(�D�%i�J�� 	���7K���e��Ė��`$yS54���kU��/�{�r�g][���>���8�UpO�4�q����7@�ɖ�;�-WZ�,}�c.�q�������l��m �I��"�������s�)� =z]:�����	"�gDi[7`����hϾ_�-�?G�N~�=��h� Nh�%;پw�f[>x��[)�����:�mO��R�U]�B��ͯ�j�h)��l|A���p��+�N��[��V��g�gF�Q� _]�X-����ˤ�)CJau��������O��D��t���-Sf�Lsa��� ��>[�p����$�Y��v�Q&�q|��}�x�IҤ����٫*(A��t�ܲ��RXM��l-�h�/	�q�!��*w����M�K���h�>���<�[xhͤt����Aݿ�<��K8��p?�E[F�(Ц�f��Q̄nD�\X���A�Jɏ��������˩Y4��œ)�l	8�^A�o�;=�v'�Vҿ��Lİ���I^�:w��Q�u�mg���s.�W���fc��Ɇ, /�2�S�⼌+�dx���e�E�&������:+/X���ӽ���^fG��DH|�疒ƫZl��W���i��$�T�A�p�m�73!F��+���*��'�&�#k�D��������&d�.S�W��4��� 6#��C�|.��Fy������9��w���U�T����X�N��c��[7�gζ�����`B���8r����	z�F�+�'-!����BLL<D��ػ��.�}�  �h�;S�gS_�e��x�<fA��r�����[m׊�r^�oz�dX-4;H2mcG�f�`�RP䥨��4��Z�d3*�8���:B�[�y%�&�%�t���)�/��~#����[d��B5ϋ��.j/ʑ���שm��Vh!�Dx_;�-�Zm຿j�&_+������6	���ge�QQ3uÄ#��ƾצ�Ic���Q��v)�T1� G��!�̱s�����Ŕh�܅bR��IQ�B��OAVg8���T8۪��d����߳�t�:��m���%z�eA���N���&�� Ȓ�%o��\�R�?Åm�1y���@�#�a������Y���*��9�B�d+��o���*X%�:��X�a BBi�%�d���7t�n�>펻��� �ƫj�a�Z:�h�A{}�d
v���Kj6w��6�?l�Say�q�e&|f����&�_=����>f��) (t�脁#<�qո�V��Y2�5.sxL�x��I�F�/T�*\y=(��mT��-����I��q�W1��zka*36��K]�f���6�(>����	����}i����;�,�������i	�Q���(�@��`9	�[Zy���yuG�Bh�,e]M����:�'�a�y��YGl�E��Nb������K�a����(�e紋2@9
��[륙p���-��V]�Q'\φB^�S�rf���8=�v��T��&/�Q���ݩp3�9��:p6kA�g�9l�D��y6�(�^��(?p��=ŹƁ�'�g>ڔ��jd"�evt�д��%��7�D]�o�$m�:�ls긳bۢ DX�CX�C)0-J��wb�9'���g��F;q���5&��Kwߢ� ���F5�M���B��Q�B����:��*�Ry���'[�Qo
�B��M2F�X�-�j�-s����SewZ���TbĂj`���t��Ve,�:M�hF��{�e��hrxM�q�T��enx�vC+���h�S�(��a���{��T.����gС��?��{��yn�=�N��� 6a�>�~g��/�MrT��W�u��A�2� ]�lY�����NpRDސ��]R2.Ȩ�"�ՌTT��a/���2UV�$�L�P���h8*(x�mj���+�;x��؊
�������뒞��#�K3�j����ל�z?�a��X��`)�ԛ�-G��t��Z?H�fc�(�Z֑�;�g���������F�l,d����I7�8؆8U�3�EE�҈:�\���-�����c��b:HӞ�`��L��ʿ��<��B���W�J#���{d������Ŏcv��G3���M+�u5�Io5���mC	'S�/�OZ�v���y~J�ړ���&A��X��ޛҮ����h�Axs,�����W��;�ۥ��*�D-x��CX�V  w���L�� 2-F�=����^c�$"#��Bh�DzZ4"7��+2���]/�d�H�`�����?�YN�:����&tv�gI��QFJ@{�|�eT�_e]]��vüa�	9R�Ы��i��rbǙ�u��r/�70�4����fCu��Q����F-�`y%O")m�ЁA��TUxEB|hN�1����͋��?�`�������[̴7��W�����`#�9 X�e[	!�g�	�t������J!ߵ�zf�;?�%�+P6��}����	|��Q4+�YT7�ulՎ��ۃ�K1���� q���ffy�r�qS�$~�LP�f����Ii�C�=��5�{[�t��Q�#MȈ��x��v��y���^SC���A�� u�~��G/)�����-�����-왑�Gͦq�}`5�z�p&�a��P�j�A`�0�XK������G�MUq�G��ʬ'��-�4ڑܞ�� s���6�ۅȱ��t���4�f���Ml���8=��7��ݽ�j�)Ҩ��q��&#�"0p�{e�AZK{m����o��A��C	�k��$F|�A�̮hw]$#�wJ�ФN^�;Zm�ga����YT:��=�*��WQ� ��u?ZqaK�}Kc�mEQ1�ڇ �\<���(����5��c �_�Z���ΩQ���U�g�(����H�,�h�](\)��E}����yއ��Pѕ����.#����U3�k�FF$,�.��0�\�fQ۵y��PI��j���8��t�[�ӗ��f���z�v:��ct�i�ԑ���1-$O,�в!+6��g��$]���.U:	_
)�/BM��^���_���j�\l����nr�X�'2L�b8�i��T�-�����B��Ĕi�r��D�>�|p�me��&[Lou�L�y��ڑ��$�?�h/P2�ya���m� 6:FP��� r�T�M���fhG:1o�K�)��ɪy�.v�R)DJ\��F*35&%v�Sq@�c�tk9���,!�.KO7s^_��ې����*Ƹ�,�7�6+��G#��۸|oN���λ����q~����I��y�O�ו����G�9�r�>���[+�������	���=�{n�VvLn������;Q	���+�����rؗ�;y��|�=#����#ʚ����V|��{W�-Pv/C�XZR�>|�[Ӓ�����S"F ���0��]p�9�.�~��Ԋ�N��1W��x�;��p;Kj�@/z��D���ä�a�4���AI�R�o�E����ΰ<,��W'W� Zq��G���}<Q�h�Bqy&ttʄ3�8���,[+؅�Hq����,Pz��q�lo�K�I1u������:�p��m�!��~�XFG���x��S1L���HkLa��v���Z�.�� ��a8�̴ɢnjXl'��&���I&���ܻ��C/c�&��W\��_�����>��X\�g|w7B�l��ف��bŚ�I�Ҍ�9�/[�p�v�0@��]�CA�����s ,�:?��T�!���:r�9���l+������Q�2}���������6�R���[�>lw9�y$R�������b?��1y��ɜ]v1[�-�O�[Y��r=��D�ƙ�8w�,	������Q��8
m+���	�p�R�XGSV�
�K�(4㔙�ˤ?4��z:����QJ�_��o� �ト�z(t,/B�%0�=��y�>*h^7	S�7�4��/�
)]ʰ�ym�Qs�w��"��vϛwB�,*�g,�v_V��H>���$3Ғ��B@���4��SN�4���{��~�ʣ��U3�� �]/8�B�M��	��E�QԐ���	�弰<�l%{Qq,y�p�f�|3h��Pħ�W�w�Mj�$�I�AF�(�v��Wr�@��Ν���1����$��g��Q�g���~�T��,t�#��D��;�%/А�c�GUY*���.{iW����fx1����gm$�Qإ�2m�UЌ���֧AӁ|�1l�4��gLL<�_-}+/��3�@�m�m/���؈ht>�s���$���$�}QH&��Ͽׇ<���K�������qo����i�"���P��X��ݡ���i10��۪�^EA5B�,�9�����Z�@f�4|��g���3`��q�5(�}���t��#��r��:�ي_�h_9k;J|�������@C��̒y7����̐��.-��8���	��v涂�5�*��+�uSڞ��N��N���r�E�fB���A�{5�@oA���$�7�C;�@���&Co�<��9߭��M5�@.o�o�#-�<=�%m@���x�WQ������@��.V@� Գ��${B��
����-��1�H+�������)� ҬҺ�a��w���;���w�����W=�V�� ��J��t�$�C%�ͣ>����✛B��3("����+}ZP�k�15A̵ɬ�M8��%���Y�6U�~��M�Ds{2�5��~
�:Pfgvg�S��8͎��~m��a��U�u
[��(0����%���w9 xM���[o�1��:�KJ@)��Æ�����j��#��^|+���n�� m���y�s�;
�1eP���[�f0�bh�C^©Wx��'	v��|{� E.�B�l�@W7�v�bYo��xs^R{*�|Z�g��k{7{XJ(���\^m9!�U!���i����4;I�jv?��9�h4�2�.� ��S�ﰰ�4\S�ݵd"�W�Y��63�&�B6�'B8���lY�֜{�L��<AX�m���N��I����1�ٺ�n�Jq�q%Z�f6��6��$@G���yfZ������ѐvD�ĕ&� *����E ���y����`�T:�Q�\O���CQ�Bª�Uܘg7���2e�@R�m�t�Ήf31���-M���űV)EsQ�\BZ������n{Ef�#�@7J����7H%���2ϭ�"|ω��. l&oa�+�;�t�{�)?k��w�g0Z�-����"un<�m�5����ɺ��K��MNr'S��9\8��Zav{������,v��H��2�
P�(4�ϐ�'nꩺ�X�bִ�Qk��(r�r:iˈ<���g�U������\ﲶ�|ʄ6�2�!��{� �*����2��?��-(�;V�����V̕�t�(y�!"�cm���p�����jT�zH����['��J���^A���\:�������/��[�������[����j_���0N����UF�X_5����ٶXK��wjl��|��(Rd` ٛն� �R�H�X�i�hNx#%&�L��h���r9[���#���K5�����r��B���+)��<O�����P�/��+�@'��N�U5$�G/���*�7&����I�^��Ju^@�݃:���4<�\��V@I��q�V��9�k��3
�RqK��=:�d��$�-��� ;
l�a�O��_�j	�`h�i't�q��������g����6�!Ѥ�_�d��l+q�9�2X:e%W��i�qΡ�0��e�����Q�")�I���[Ϥѵ?����O����{��K�
 #�T���Ч��D�~Z�g)�f���,`��@xbϳ2M%�k�s��Yrĭi_��ث���{*I�K~E��ʍ�7���`(�%M�?�����S��Z_�o]�;A��A��v��S��e��d�� � k@���=U(|ήs�٭+$�3n�.A�����%�lI1"��nf�`$Iy�;�ޜँlYA��xw��I_��[Ҝ�;��x��(��J��ѹ�'v�J.��<��Krd2�K؃r������������Jʎ�����{^��mP��뜎�xݣ�&��ɿ��� �q�5M�ynI��� ��D�.���:�Լɾ�2Ϭ��;��H8_�j��$7��>=i�֐���ba�g(�g�,7CK��V�we�C���r�4�����B��ܰ�u�(��)zZ�:��r�ECE���(���+��?�Yk��� ��N��4ӎ����&�Ρ�nWku'=�7��`��IE[��+�x�&�%sx?�;�o=��C�W�����Sn�۔~&>�8̿���N�6bK��&��	����9fux��h2�3�]������Y�!�o��'+�`GF��-<�]�̖�*2"g&'��F�ˁ�4��g�nT[A���\�E�of��������f�Iy_�d϶ӭ� y�K\!��9��MO-��V�Cڐ���%�� ����f^I�ȡTT�H1���-��������v��	1_�D�9}�ԔK?�SG��gÓ<ʕ9 �R���^`�Bv��Q!�/�f^I6e0f���&Xy�F���DgY2��O�i9mzI<�"D$}#/�����~|.CC�SxϬ_�tK��:������$5�V(?]Jaߦ�-y��p��*UWȿ�Q��Eڦ���T�n�n�u� ^0鄄2�e�w�@�~rm@�\�]�E(t���4ۗ��4��`_)8�
�\Z�RO��<l)�ӑ]0@�@߱�]gw�\V����R��{��M!�ǭq��{iC�-~V�t����$c~����l�k��	?���_�#q�fk�qD�k�$'�\�|v�`|B)�Y1$:��l��U%��j�a���5I>h<a��A��P�	|x�7h��^W��K�8җɌW/��$/�ؼ��!��6����� ��A��Pl��^l�2vh0�ڝ�ʎO��DO�w��lq��­먷�0�;v0��FZh�o�c�₡�˶E{�b�(�� ��h��3�7Di)#dZF�۶^n�3\T�4詥�Ls`M��#�Y��*"�`��9 Y5_V��m���fQ� ݁<%�ĥL4Դ~�k�<��tN�Ubw��&��:��b	��p%I +��$c$.w�sZ*݆H�%�k�>����f��Mq;�n�%�`�][�8��*k���Bn�S��U�T,�wx��ؕg�X��/~�i˂���kaD��h	m�"�ԥ/���K��#�����`���MȒV������9�:N� ;��$���0{\��B +�RDޔ?�<�Z?�`J�
�Ƽ/���a�(�ࣾ]3����	>�3��x?��Զ5�D��ljlˊ�.�*�u�)u	R=QTV.�g���v�ϖss��N~����M���/=rr�ta4������#5���Z�ʹ"�,Fʽ����Y&T����D�6��p���V�r	Y��x��7�����Sʕo#��i����|��Em}?�ҢX����))��o���t�?��(M�����k'*�B0u�*`�``�1Q���+�3�0$�@����7nv@�ȭ��i�$TF�x���3e@K���9`��Vw�����(\9il�|�5B,�Q����{|�h�q�]z�>�~�A&���:������4R���F�y'n���S�H��D����L�Jv}� ��1��l������2����G~g�q�&�f�6�%�a�A%��kƢa� S��T��w`巺`�f����1�\q#��z������c����d�\
��hl��U�>Mb�w����k[��I+nTQ:�E"��5�c�����?˾93�oǬt�'���0C�G4Րƫ�CIP�� Q@���Â%�`Q���jz����u��&V�W1Pܭ�C��l�P�Z�5�S��+�U�aףk�0g���"��1���o�bA۩���?{"��(A�kܒܡ�#��g&i�b��S?a[�
���-W�	Sڲ��B���Ak`�W�郐r)����	i�/YVo~��@.xt��A��3H�!��[�EmAq� =�d+�ֵG�x0��� �I<'����7�vD�ʵ�W��¼0}5�������
���t��u6�(z�?������!%�������H&�Yjs�U>C������D�1�DAY�t(k[(�����_�̮r�'�R{N�}����`��"���_O9g��O<�ǘ��/�u�d���>�5cǊP�B�2�k�����G#��;��NԼ��Ќ֍_>�	Xg�u�AcD�(X67��0�J��@ub�J�t�����M�K �`�>ˍ��4�-�-���O7�.�R�(8Q�a�ij���╚���,�超4�%c
�9=����4t��'`
����RqK&!��ә+�-5��{��q��am	>z�T���ʝ�^а�·�?	MB���efب?UU?�w7�yVy��$����+�GtY��0 ��V3���v&o�^;忳l���}ʀǻ�g>FP������gE06�\��*���ҟ$��8����.������M%ۥ�]U���+��P*~�M�{���1�G/��͌I0�/�n� �\�g�A��͍�k�r�����4��=�v$�L�6�^߷�Lmә�8��8x%� �̹6�����,nj��zJ绫��g;W��B�u<�v����hqw���NK �3�c��&���9	 䃝��Ti2�z�D�������[Q�Z��92�Gj�Ç�8O3���8�5�R翐�(2�|�r�J9�+i�o�萺��z��J���=�������OP��~�p��X"�ݗ�ƛ�șl8�� �X����@��Y���ѕ���l��&��k�M��'�|`9�'q#�E@����� aQ�뷦�(fL�'�ԋU-��N��E=����f�{Ȏ�Y%%\��J%w�`4��|M���;#��e0�̋���;���I5&�)�?���敱�R�a��S~'�Ҫ�EI���ّ�V�f�~��ӽ]���3J��>�
<
�I�Ud�jL|�ҧGd�u_��fa���9�Ff+G�u"�D���/	�(�\�2����]�,�;�����KF?��+%���Gל��l߈:��G��q	����B;]���Ο�1���(�|�GB��bP]�s;>��CqXef��T���ໝ 0�c�YcW�ؠ	'�	Vx�<)3���Ƨ	��1�ĕNy��{ �Dۈ�gl����
�㑬f��i!�Z.ƍ���v�ċ�a���}�g���w1��� �R������, ^�[��I�+�N9f��?���d长#	m�j��3v6WQ�5�{G�����ng��M�'i�ƨu�2P;��.��6�r�)���HX�!c�!Z�ezt����]�$��|󫩀��"�yH��)��FM%M�L��鶁[�c���}T��lW�(j����n�G�U�B �$8K[P^�$��c.Ka�ڡ�	<AJ�Z�PO�X�|%�	z0�͗��҉<�̢�Ԁ��<ٷ���c�8�Z�*P��������4��~��̲�D�`B ,����s	t�L<�ҷQ���C�Rd�����(��l�������um;p��R
��O}Ӕ��Pf0E��o�$VJ�����ho��6�((���Z�*�U`}��xզ�K3��!C�s�g����R0�L������YݤT�y]� ��T�(dV�tŬ!g��#��Vf�j�D��`�z�X�Fg���[��uo\���Xs�T'�������N^z����	Z?�q��K�	 /���M�C��E���ݓ��	׊$w�ӌ6䍋�6���1�ir\�z�C�=��&�ɏV��}};f��3�E�Qq�{�}h�:}�"�&���O]�|�n
[����F�J��0���ُ�RkX2%?��Ūm-�-����=!��S�G�c�&����>ԩ��E���o=ӷC����]C� ��F��Pi��T�Jbd'loI��\9�v�@��6)�@�%��:I��E��8F�.�Ѩ+@�+,e8a�؋�[t���������6]�R�XA�^���:�L�͝���'m�G�4\��{�T��q�}s�	�x]`��*a�y.�c��9w�i����	��t ��bǌ15�e������k��(�}C
Y����9�|�Oֻ@�ͅQs��9�à��=U����OQ�Sb{�:� 0���T��n��gLW<��ЦAT��O�#�C,ؙ�Vƽ �[�V��������1A��P�H���v�
��\��ƍ�@r��TЛ7��s��O*HQ�'ik��>���N��Ο(�@m�{�w9�,x�����F��p�)T���-��T�E��i��y�������;|������x��8ߪ���V-�MegCd��j=�p�W.Ǿ�MG�K'F4��z�иf��m�~pIr9�v�+O2�\M�榊)�dWôF�/��漇�9_/Vi�j0]ٱ����O����RXǬ(6`�!�#F�uk{t�a#��;d��tڗ�'Z-jMQUdSm��nY���m��5���#�$�l��ʤ��_��k��_
COf����ۊ��G4�$��?�3��v�������3�
�T-}�L%Y����������H����Ґه���O��-m��0�'���_�6��~�|r�
u��x����x��}�`���:C�o�/o�z�	ˠ��N�a�TA�z�/.���*�X=\���P��W^�^o��Xi4!��C��l�?�Y�����l��. ~������~>�Ͱ5�¢m�TF�·F��b��L�Ym�5S*���E�3=tm
��[i<��P�e`����1��8�o�LZ��qU�,��U�ʘ)�WX�Z��FU�
v}��I�c��!3�ۂ�0��O�"+���Wν9����Y�ۆ��j�$��ϋ�.�'�@@�F��Y߉�_�&�H���qI9���{ʺ)N,�NKp���=ck�@�p�TY���eʉ�R}���l:9��i�(�E��Z����F4B�DS�g�^������x�Df��Y�SҸ�i��
_2�=2�)�4��k� ���jœYo'��4��!��J1=��҇˪���*m8<���&�@���	�6m���%�K���9��Ǧ �E	��orD�2���ġ�� ���̟�bAQ�
���>�.n�I��M[�c�7�n��?�ڛ�ܨX�&��#,p��W�L���).�A��~<��%8�LЉ��}0��m#+���U.��VP �Eq70JR�Sܛ��^���#蠎������E���(1\����?�LFʏ8�f��}��RV�|��e�u9��͘�R��%�����MZX���ݐ�4w�KC@W�ܨ����l`�U"����*���t|�;fm�c���yu�x���	1���ک���zp
���֔�ݽ���L�`	w���]��Q��8A����f_U�5���8���v?��V�h(n�6lQ��H�AKc.ˁ������9�,��N�D�h����=	�B@�a���7��4�W�kN7��(�a�HN�ȀD��E�D�Hឱr�p��/�;20�Ex72&5#��@E/�����5cd�r�`���-m2o|��vi]6�z㴹_kⶃ��Ti�4��a�P�mCCpr	5JԼB#���@�L��U�=��e5��O����E"���0]�DO��S����W/�C��������+���e�'�p�f
�y#;��E%��~��gS��$oaMN� �o�i�t����ѡ3��� 9�2�2��#}�)"n�R٤����\�A �����	pΦt�"̶X�s����p ����i@Vb!�̍��ո2ֹ��q�ɉ�!u�63q�F����%�!<\\I*���D����S�9�SMW�Pme7���G�\�d ����`�{��Ϫ%/��3�Q��$��I����U�Ų5b�}���j�A��z	��E'�v�������e�,h��_���ƪp��E��P6��`�L,�uFח*V�*!��=��Y���z#�g,��~�:�Ɨ�����M�wR*_|�*!C��iFo�h��|%����^*�M�H��Ĝ_�V���lr����!h��¦=�7��>[ ��x �u]�	��VF��y�;�������K6�Ǡ�}dZ�O>VF���1��Z�a�H']���7���
�e�2�;��3&,�����Ӯ�!�%U1�襕��S�h	`ws_��":���z����S�@b�	��,�����G�F�E�d�8hD�BV���4�[G.:��q��q=�U�_+q��+�C�AW{�� ��\Q�3C՗�YOǹ�y���Ʌ����|���ydV���N��q{j�}�� �O*%���){��+~��
T��wNd��`ƋA�z,�@j �e������Ju�`rJ��*xl�L�����7&4i�N�<\b�vC��kC��ɐ+EĹ���!b
�'w�����ԩ[�Aܗ	,ŵ@;�9���-^_���VN r%��!�L[
mb�pRB?7�+�k�W�s�^˚K��$~�g)�Ҟ� #ab:�^@�,�$��Wh!���hO��@�6Q�q�pՁ��J�Dv� �7������:�9�$�Ԋ��S����2�q�Y�i�2�l+�`B�%)g�%ǉ�T�ne!EF	a�[�އ�1$6�<����ך
~�j�S�VJ���Q��t�_+�<��Śvv��B�>SV�����Be���R�J����[�ʏ���B*�����)�O~�&H�*y#�*��_�ږ(~����@�I��M0(h~���d۳�����Qr�^!���9��NU>D V�r%k^�0)R~�]�%�AY2�Z�$��-��z�-%�gX\ �]�GC��h����c��>���JV+�ϡewZzL\�e�@��Ȅ�y=�c@ЖT����FI�~���;�i�9F:�1���9�_}f�h�8�nv�؆�_Ќg� ?WG�x��?�I^:�� ��Veob7����'��8t]ש��9�@g��PI����r�@o)D���4��⇨J��n!�m.i�PS!���Ee�	��	u��K ~{���}Q��u��#:eY�`�*��M�K���ϼ<�6�#�׈��K���8ka"Ζ#�E�N�����6�=�L��5� u!�n���0X窱DbkFK����L�g�v��ݸ�	�*b�m�Χ�]��e��:$&����KP.A�:����K�~L�B���gӁ�f��rng��_ڄ��(��>�w���1M�Q�X��S����Sm���>��֘bH������� 9"V��ǰ�6�~�S�*2�g������Jz<�N���Qg����7��V�n'B�͈�Iu�����M��<!bq���n���sg���]�B"�q/�����0��	;�=�2����[v���|��Xw�9���j��C�$0����ذ2ԍ*/@|�gRS������/�>����
8��$�@�l<A��O5"'�b�{f��s�/�-A��k!T-2�ǈċ�I	���0މ�*A�'*��#[�:����Vq7�%����!�@���S�$����Q׈m�;�ֺ���F�7�f�&T7o���a�F���mn��A 䳔��kz�h˞:�?p�/����ɮernD��ؖWx$�H-���]w�oY���0z���DPGR,�ߝ��Y/���C���䙏��NZ�\�Ke�S{)�u�w�"�v���R�Ϥ����
$��R9�v�I&a�BG�� ��kB��6RP �b��S��P�(�PG5������W�&�(CW�����f�vҶ�ęޱQ,g��"� dSI]�O
�D�D,��ޛl/>����e�:omԭ��b�p� ���j"�F*?g�n�~xE���.��Ik�9����qi�ں��3Ml��sn�ɇy�TRu��U�ʶ����}�v	)A��=�ų����z���� Hz"i�M#�v�'�; ����S���7izE�5��r������K���E�KW�OF�<|������ʭR�� A �B�c�L������@��<m�m��P���*j����]����-z�׃�j
[.o��@���D7a�&�jc^zҘ��5,�D�.��ԨZW�������|O��������𞁳)�P6�y��EĿQ�<B���o�Y)�4E�BCDb{y�JLeA$J�&0@�:���X���hjfF*�)����]�P�Q��T�d+�}2-P�kg�*��ɽ.��U'�k��d����ٝ�,:�0x���ߕ��}�k�\W�O�y�S�o�b:1rď�H�*������s����#ܩ��4�8F�޶��,s��+�ς�w�������˨��YW){$��W��G�O����sUD�����nq�S,Q��S�����gEݻo��FYe��/"�GI��|�AB��"�K[�DsT�?Z��7�^%b�ä>��+aΔ��	�S
���8����a���������P�����㳙�~�A���B%��mH�۾���Z!{&���I����m�_���pg�E����NR�gg\&VKIW����z��l�|��7�7>�g-�7�MٙJ3��7����HG�B��ȿ'�K�ҫ4 �
˃�4�8',�Rc�>���m{�������w�2�=w�=������/�Yn��asD�����4��_�r|*��u��bյ
�Y;v�T��.1��Z�S�ƓŒ8(��4+#ٙ�ݍ=�����G��$���\�M�=j�I�N,��bS�J^o`�y$1Zt*۱fƂ�8|�kP6��+�#3Q����.Fȥ��B��S/�Ig��fj��6:`d�n۲�l]\��(A�^��_�}5̆�d^=�T�0�=����e����#�P�u���~�ʡƉ޷�ѡ�J#� �n�VJԾ� �'�	��m���e�Ao��kb�X�.����a��(:�\uk������-�E�狺���Ж�xآ=��2l���Q#U-�nA�5�¤*�S��~|�P��)�U�4���E�Lj>���F�-�[L��p���x��2�F0�6M)_�� ��:;-6�E}*��g���#�v?U��l�H;���c��t�JM�?_ ���.��.����Ơ_��lCe�٩��Ч;��z��T���ow�����@CG�y�]/l���&Du��ILsk2� *A�k�l`�ʁye=��
Rv��"0��zP� �FW�me�v��\%������ҷn�<�{Y�# ����J� R�vE&�0�!t)Ȫ�ͫ%�laK[~dN�{��Z1V�g̏����WYh�RE�B�n32(�0Q{���W��H�ƽ�hW^/��R�oe����+�֨�k]".��r-'+�յbѯC-T�$s�jf���`
d@�|�q�<�H�rP��M<͞7�__���Dߨ��zY�Vq]���?V|���gz~";���[���:xY��_�Q Y��d!"(5��Z�>�Xz��[�K�a�r[����Z>1u-�&�߀��)&��{\��,� W�e'`=��f��%в'pDV�N"����tC���S�h#jn�j��p��c�U��M���~2�<��<f2��Y��+����S<�م6��	s�6#�yqC|��
��yD �]Vğ	A2J���ж}��?�4p�(��(�8�Tھ�E�����t�l��'����G���r�A�N�'bɐV	�Ŗ�� �b:��U�K$r�����R���{ ��IIA�{������������4�+�A�Z���q�&|VۂRIF�/��f&�[�B���\_�Snw���wD	Ԇ���ս{�Zն�pL���M6FɅ![SA&w�I,"�U�ĔԆ��̓2��sDγg˽���5!�1�ǚ�������gt���p��1��X_<43u��R���Ƃ�4��Cs�����ٓ