��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&��n?��1ů��> K��D���yE�42i�0 5��l�R����꨹<ڛ�\ �*�L���T���DL��3S&�dC{��$�d���T-(8�n�2����L�*��1�8�PJ&P:D:c���*(�w�]���4�x���J-�h�ҁ�`�щz� ŉ��Õ8n<�1$կ�����鰱� 3Z=�e�7�cK��K��F�DE{�!�v�:�":l��:�b;?%�}�5���p��yH�,��*�h<��p�)Q�C��>��=�?����} q���T�Q=Q2^��0Q��P��'��t�R<�k7�6��F±|�Jb-j��Ǻی��r���}��
�)���Y�`_�A�kY�{��>/Y6�
��u�4A�j���ĲN�ޘk�V	W����ݫ��[W��
!0���b��p-X����aF+DL��+��R�(#:ڋ�����Z���v"�9�������BK�f�d�l�2A΅�z��-搾��,��O���NqK#+j�W$=r�J�ݎ��c���25q(�Ld�$^�F5�O5]nc���e6u���6ի݉��˛�����'/���y��a�nB��	Z_��t\�X�� 3Vu�G�s�7w�{/�)�"���]�<����([#�x�/��>�%vr-P]��p*�6 .:'ɕ�D�o�Z����&�P�b�,~�v��f}Oũ1��T�2x�4��:���t[��[UP�؉����ʓs�M�S�K+�Z5��`�+�Mm�I����D�G��C{/ɀh{OWߜx��V�v$�GN�Џ	�U�(��*�#�NS��n�!P�
�Pdw;��X�1@W9�È�ݓb�r���I/� 4���Ë�}�0�OJ����"J�ut�S;F/19�����Օ")e�0�'U����}h��[�����n�2�{��|���yJ-�J���p# ���r��Y��i�a4�_5^Yy-��e-�}�W���_�ߟ'C)�k�E��Y���������?IGa6C]L�k d�C����2�TJB�^��)�A�Ԩ��z�����X�t�	�gV� ؗk�R@�?��C�*B����	�U�L�����D�3Q�����g��?l����3c��0Ԯ\d,b��4�,��͟��DMG~�#�[gZҫ�$O�`1KHԈ��O�3�ʙ���BY��w�Y��f=���q����D�LЪb�rmHWl�t���}�& ��҂åS�
33���'mڗ��GM���eq5m��ND%���M�m�M�{!D�D�+�h�vK��w|�v���U;�)T�hޒE�~�? �y���o�]-�z�A~�!�u�<��͏h������Q�#�XgQ�Zw��1�fm��x��������<���-��[��>p륳�z�A]6�Da�xl2+������>bu�3�Dwjb���ꞟ����(��z�{�4�8+U�"?�6='��I���ڤ��+u���S��c�|MTık�_+L?|$�7���{��6ls�ݔ�s���?�ͧ��)Ŏ�:MCm.d*]��� �:�;�`��T푷�e�/A3�	و�A�D�|E7����C|�O���%6o1/ףjj`��n�31�2coq��cp��%�xx�M�id
��Xpv5S��T�u�˫�8��Z�[%O�3)%/����a�<�3�z>����GZ˘���bt�t}�8��*M�(F.��b�e�d7|>u���K�H���C�jl�C��$�~r���Dn����c�9�ne�)԰��b���Ǩ�52ҼCMcI��V���A:�o�<?�����}y���/]�
6,�S��	�+I���j�N7r���ϱ�������q��-����hs���d���t֖Z�>Ő�D4+};�h��n��Q
J;׫g���@��D�!�����`�ty�yy!�S����H����WUϔu�	��0S5����C��1��;���?A�F�)�M�H�b'?6 J�ǳ�^kyAZ�G�z�6D��}殊�!�va�7�����@PUuV*A6&v��W
���v����?)`$��[+�0�+%�"�@�4��ee����za����<��	~�I�O1e����a���f*?5��X�0M����L��������XV�ǥXЯ-R��櫓x�#���;�ԍo�J�����&��y6���w{�f����~�=|��rE��[�Y�*r�#7	�#
���K��}�Ԫ|��F��;(�-Ӡ�<�j��=+F�UV6�~�F��;�׿�A��ш�gJ^2R-�ݫ�4�+68%	$k�	�	�����VhPo4�a��T�ӣ9�Q��vxS��|�~�ӥ(X��
=��.=�A�݇�ɩ�3�]:���KL"��n�dX�[���A����?�N���,΁4�xډ>{�̳�o��	��^��0�����
��O($&f=x�Wgk�P�lk,m�4��!�����`��ɴt���0��q��̕jI��Q&#���d\D�X}������@�W5!��ҟ���c*i�d�:�,)��aTUo����a����,~p{D����;��E�7/jWL�v���S_s�zW�.� 厣���ͦM�N;I��2@�kt��p+��7�*�Ût?+�䧨oy�ȋ��e�)U2�ΐ�3q���*�S�]O��T��9!����D���a����ԣ/���C���^��)�q��z�ǭ��Qt�x�Ĩ9�6%����I;ќm"�W��@�ދ��Tp��f7z���9�֠X�3̐��w���W˹�f��Aq�t�?1Rb��Y@�P�`\�x�o�K���?�� s:e����,y�
�D��TB_0�@�F�P�/(Jͤ����S��#�Ԑ	lʜQ���#tI�ׇ�K)nv*(ySȹ�����bb!dy!0�����b�"U�h�j	�'"�"��U.Ir�!٨�t�*v����"�ɈJ�OѢ��&J��HO��ph�g%�Z��yn��3ͦ���,@�>�[؊����@� ���{͸G���$���nb���^�?9zr�+�]�<O���7+�tR��Fğ 8�Ta۲r�#�ƳB����J��.��^P:��Q�RF��w?xB?��m_3��BĖT��;]B�mp�����H؞����Z��Q��/_U\'��j3>uW�ƳYBI��v��}/�WۭD�5o��`�/�DjMe�����LU��6����n�8㲚�(~��z�0�W�+��e��3��f27q,���S�q��#���͌�r-��B	^fc��4�����b�x���������,K�P1��xN�R{i�⽷���sE����i�)̓�������e޾ Na24c/����H�P���������W75�6������+2W+k�WxhU��j�����2x6����`
�(�&�t�`$ �:up��X%���
.�h�W��&����I�����D�K5��U�5��L��ܦ�
T܃����5`r�s�Az���em��=&#��DK�@H*4���;����[�تF�cf�#]�mL����!�8�j-���\t��?���*��n�*�$ށ(����������e���W1���f�Ԭ��d��r t�J �����Զ)�N!c�Y����I�}�:Qǝ+�'�n&���
�u��&�� "�+��j�t��'S�['׍'��J�e���c#G��r_c��[n��A�	����`���fB�O���Ȥ�h�7I&�֭����X� ��AC�Q5L>|M����z�������S�MK��-b�v�.ti	��Az[�ţ���*c��c��F�,������K
��ťF_j���M�,�K�=�z~�ʰ�ód2xz0`+�����İ���b�T�uh	gD�ww�}��:���ʱ�� �YzeE]�9�t;)�4��j����?�I�9G�����9��j��'������~2,W��ɩW��U�h��|烇��K��cDh�7��4�Z�姭�����х#� ��9Ϯf���h��Y?%qPi��w�"^F%��Ƨ���`*���:�N4e��ջħ��/��Y�]��	�Sb�tF��r��1�U�Q�`���ì���hZN�Wki�F#��p�8Ҏ� �0�=�=Q��c�fl%�]��L�NWNw7��U�sx2���.���d?	48��(D_M���o������Q��8�6��S*sdmtc�Aq{Q���1�G=��b�]�#G(��p�b$ٝ*jI�ﲯ�`����U�!_+�)<k���i�ڟ����4�o�͓�7W�+l�Ӧ7ve�Fp�Ts=iі�I��3e�T��64w�٠����r�&4;A�j�炌3	�o�7�K�ò�zt�Ͼ�^S�^���A�{X\Jl��8y��̎R�|�@\=����󅒷����S������߄�?����,H��XP��/>�֒�i�ҺO<�,�Y�f`G�p�ő���ԧoO>)qF�Z~�$3W�PO*�Z+�+�d-@�
�k���Ȇ�R��*ǡ3=�21�f��*�r�gǍ��
�1��˃���Z��u�;��"��{SwD�r(�u�k�0���!�۝�=*���
[�E52R�47N�ɒ-gt1��,�����Q�]ήo��L����;^ ���:rn8�S)�,�;���J���8b$����X�,%c�Eﹼ���g?�ٱy�ǧ��?'`�/��A�-���0�@\A��oY�%h�r��"�3���V˺�@��Tn������G	�q�J�� 2�r��H|��p�fV7[�hX�^�q�ӽ��s���#��	�E\�@���/����a%=�ޠAN������6P��7f4�����k����?t���7j ��v��?i?'�Kf���^�/�6a�h�\�����O��|�=k��>���"�X<�S�ƪ��ۏ���#$Y#�ن���|$�\[����@��'�!Y9h`Z��z��O@�Pl�T��0<�,u7���]���U�ql�DL<nKK����WR�vq����ܵ�r�
�C�~4+����Cn8�rEA��M�@;�+Õ|yՎM$�f�u���D9[Yf�SpSA&��<�;���ɬg
V�:�W�j�[�zp` Ffz�2N�B�������)[)�O�[�GM��`�6��9�+^	���V�(m�miH���̈́�({)���4w=]:��������*0�z�m��Q7�.{D
�1��(����
�)uw�<K=��UL�e0� �BS����C�lN�>��~��D�-�5rV��Ұ�Ji��/��/�"<t�T�=&��{=і! 1{Eoǌ�M�J�| �P���%5r>�\����n��≃�gLpГ��7��٨hg	ߑe�ϲ,�:�O=ۿ�&o����o}i�T��(�.I��Wq����l�k/�x�&ס�*����Fz�13���ي��0�^>�'�mJ`��LM��ƅ~jh������j��~���C��U�2Y��j!��R��vn�#���q�y{�nn���� Y��-/��,�
u���Z���=�y*�`�t�����9m(�Ѧs]U�i<-����r��p�W��A}�K������T�p�'\ MZR��tڀ�xؑ`F@����2.s�r���_?�$���b3���>?��� sH`�=l�X$�'� ��)4���y��S�A�CFsmRp�8�
�;5�ӺFc �t�
Xg/���݋܏P��@�c����a|��a����ظ/���T��|�4{}�t���S��r�x�`��`���k؁�KϚEp��ҚW�~]�+i�}%�Y&����\�-𾀿���9q/��IV��w��Mmjʯ��=�,q�By���mf�h\� ���Q̢�H�`(�ʱ@q��V~Rk�^B�^$�\��\%gy$�Y	?�	#X1�E�CP��`p⟘"X.׼&�Ԥ�0P�6ȊF���I2�i�~va�~����� �β�T��Lj�<X��ti���h�3J���O������Hu�����2s�h�;��~���u��:�3I�Іt�e�*�JM�4��� F��s���J�٥.��`'��������4uNI��f\Њ��ݸD=�L�=��"%[�� �7SF[��B��`T߇�+p	�񹰓�꿥��r��|���I��ꜧ��ҽ�O�z�0��g��D�m߇�8���fj}.���Du�� ¦J*Q��t�h�jP�~�K 9j�M8�3���"�������N�)5���������]	���P]�r��\���w��s޶#R�߀��=u'�.�
3���w��9�:lR���N��$��%�$0�l�?9��7Eza��3�E'�\��������W��7S��
B�H�����H�:$����5sə���~�7!�L���w]퉁�q���f	:I�煗�	I�
�x����b���y{/�/�Ֆ��u�c+J�J�� B�]���W@��\����v�!�|�i�Fr�9�g�P�X�@� �/���T���zwV����:�j��<`芛�C���{�-i�[�~t5�P��rv��>��&wF�����R�҈ڀ���TXA�Y_�M���3\�dl����~VMuB&E0(�p�m���3g陑R2'��5��V�$g��	�J��;џ��
w��4uj#�8@mV��1{���**�`���8�Ƭ2���^K$	�}ܵ
���#����j���y>Mg��� �z*nj�a���U&�n�'��m<��좙x�y �i���b�+�M�`Z|�������_��#;v�`����(XvK��1`g����؁&}��0�\���"_��'���	�1g��݃3����Y�ڮŔ��>��*�=CQ8gϺ��s��n��SZ����bT��o��,��4�B%��P63͊�����%炮�n������>��*���S�S�D�.J������y��/7$s"�b�{�^�O���(���2�j��}˪s �l]�`�� ���F{��[8���=T�s��:���cT�4�Q,������U�}(S<��p�=U���v���O��23�����DE
m�������#�O�A$�!��+y=<�5�|k�o�9�P��@}H�Z3�`��+���>~*�G���ƲO+��'O��n �`O��W�_~�,;�[����r`Iy�v�]ymQ��h�P?9��)��%�����
�,�%�R���WdF���_��0RL��t��E��Gm��"�O����K���я�TH^.|0;v*P�_�0Ǻ�Q+m��?P:�����3a���y^<������d��Yp��jE�}���kB��t4a=V�9�ml�]5y:(+��c0Vz�c��	�_c�讀s^0������m�[��a�>L�QO�@������"�Q�``��ߗ4�  �����5��t��3��CuX)�.y02Il���us��	1'�Z������O��Zm�jt�Q�z,�*�ÌӅ��k�/����'��XQ��$*�%,ۙԘ�g��FH��O�����iVī����(20�>#�Tȥˬ�'����2���4ck�!M�8�BO+�~==�^�c����Ts-���=�nF�N�nS��.�M�Bk� � !�>�����%���l��u7wڈ�;D��+.��c�����$�r=�5�5e^�-��4�w�<?���(��0��R�B��ё%b�]�!z�������1i;�as��;`��,�bEW
5D��|�ύ�$B�9���k)�ˬ�Dg~aWe%�C��S������y>}fo�Igv4�C���(Dj�WZp?�|���X�H�!$6�NKxz\�t��E���K"7��m�&�X���)E���-�.d���g��lLA����e�ܥ,�֌|K����hQ�I�Ϗ��<t 	N"�+�:8�V������l�c��d[1*m	S�U���	?#��ԝ�:O��\dпT��m�l)�ch��s�d�����%82���n�8��(������PC$�?��=�O��t`-�����������u=`'����lfb*7������z��f#E�H?#a`�>�Z�B}��mE$o�?���t�3�~�7�Di܇yƒ(a���F���lʮ�7/�?N��oQ��؍���I�c�Om�?�w��{=Q#��4]h.���\�^].�Ⱥ�դ
e��l�n���T<y�})���Af�f��!�C�GY=q�/:-��3�m��c�V^� ۭ��Mq�f#slB��� ò��Z�/T�sX�چ0�	.��&o]�(2�m��Gx���*_J�b��oB<��v�G�r��{����n�B�:���y�H���+��q�\;!��L�)�%@�����ѿ���N.�O�驉��ݶ2�z;�uO*�Le$�&C^��G#�7=*vnW�a����wI7�]bC/P	�����y���������F�ˬ�b
���S}��������9�ˀ�,0
�k�<z�8�~bϲU9��Ɯ�y>�~�1Î�? �F5�e����go8~֏,�������su+w��oJJ��A\r����#���o�(i�FX�7�ǃ�ħ"��tr��+�l�I���>3��-���[��/h���y�� ����03�&�i��l5ݳ�ʔ.����3ٵ��)���M&��D2��h��p���� Jv�_�pyĺyw�k�NK)?7d�^�m����?q��;sx#=4	,,9Ѻm׏�G"�P�>�K\{E���Y��88:^�8e}�49�oC�
���*a��*"w:���6�4C}g��ߎ,� ��V�>,b�coJ�z�����q��(s��|z&1��6%��S!E�6u��.�	��g��~w�;��1_�Y|�\t~A)o�+�,��C��<&^'�Γ:�k���p�J�89��4R��wr��EF�,�h[c6G
�l�Xr;Ã��;��T/[H;q�Lr�����K>ʠ�Sĸ@���:ڇ�60����m�򙉻S�Ǒ�C���XO�ǀ�����_�˘J.W>�^�]�=��Uov5R��?��0?giEۙ�}M{�5Kip���ӗx\N�Ҝ��Y^�?�_������*�l�P]��-A��oD��|�JI7���Vx�pB��
�JSw�]�*�j�EuL��y��1;D-��(����W����A[|�k��'�;M��>�t���T�Pw oC��K�X���#��˨��5��M\ZU��"�N��r%-!����AO�bfv\������oo0�7������ݳ��+lO�����7�`i�Za���(\i2F�#6�?��(��~���h>:R~�}H9Z�����%=6D)Bf�J�Ei[*R��W����!�D����pA��u�5��W\��k��t���b��E�S8����~XQr��������yi=O�y�9�uǗ�.'�0��w�0Y�P�OO�0�O���N0� ��t��.um��'����q5����Rn��x�P��WU�Co�Dm���DT����>���t�c�R(�m�|�H�37��6`�TE��
�����Ex?�y��H ���)~�F\ԵI���z�������s{�7��`��ڛR ���C!C{��q�4J�1���+>��C����r��:���ժ*wPq�eD�+��a��C��E�L�x�*��� V�2\�
t&4A�b;�\-.Α1�qp�Ҟ�漢 �ԅ��fID�9������Ym��z$�Ȳ&���K�F�]�
�S�)6�j��G!c�l@&V�Mg����<�}��Lma��v�z������O�/�~���)G7��!�-P�4�v��W��<�8��Ó��o\z���%#��5o,���y����E��q�ؗyћ�B d� D�l�˔̈́7�����K�I�ں�Cl/�vgEB��$��R2��@/�Ì����Oq@|+6?�?%X���dH�3���.�;�h6�tX�n���;��F��S�>?-e�>��|�f�UdT��r����k� 2�
�"A����-�%�j Ձ9V���|Z��������꽂'�B�X��� ��x+�3U��ʽ��ن�u^��P2�o���#�O����Y"�=��*������I(�t'���,s(|gV�n������%hx�D�0i�<�P��v��mW�k&�[�Ly\��XF7�q��|k �)���ؘ������=��m]ѭm孇 E�z
�e��Š���&� �t��5�G�F�H�4a���r�[��Z:% ��'sc��LB���������㺕�&Ը�G��&���? Q	Ҝ�l0D�m~!�y�W;|0�� ?y���������	�d%�u�gS�;�O�|�{R/��WW�`d��ur�C��KU�l�(�a�����$�uQDa�E6�	7��95!�4���:f�v̓�o�"Hu���X
�W!�AaS��0�^Qۥ雷ӫ�\�=5N��������T��|�ڡ�^�� P��,rB	t<+72:�X��/\<�Cm%m����I��8w�)�����SfX�S�f��_`[�@k:7����>����!�j✼�oX�F���+vӈ���Q��U�Hл<������)0���Gѯc+_�A�+#NM�3΀n��u���Q���-7"�Z��T�
�
��n�L�M>��