��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&��n?��1ů��> K�-� �&�T�Ek/ֆ�\�놭5�DꢘP���+L+X�4��J��#�0�8���������l��jT��+�(���������6�MC!D�;�m�퓊D@v_p��䙋ⲝ��C_�6�Ռ��#�� ���	RD�4D��畓7���vn�H���0���fX����4 �CS�C`{��;�L����li��� y+����FD�p"��]���y��R��K�({� .؜M�������	^5���ɋ��&���&�@*���
e�� �t+���
_6��O<��7f�M��u���m(MrN����z�jL���@T`��M3��c�uQ�Y���%�dD���,�~^���y@Ga��(����C����	��G�86�S$��ɳT�ز8���:r��/y�[ݦڍ#A�����i�&<nU��<[5)�Z�-Ĭv���0t���d���"_���:�'-��d��*��q����_d�y�N-��~";#��������Y��؆���	6ZJnԷW��έ$Y�K�?�4���L�w�Wmiɶ��Y�?jx#*�i���F�m�E����O6T>]i�_�9;�!(��kH7�OS��_��[-M�((��lO�s�$�g�x7`��ZV�E���F��,9�j	@���]}<�ahb5~ãdl&I^�	v����-�@�@���	��!��d��`j[Q��� r��;f�i�.�m+UH7��/OV��c��������l��i��M��*'��?���G� SK�M��H?�ç��q;��)��Rȩ�"@���r��Ml>8!�S��L��EgeH]�8��>]GR=&���C��i�Za�z�,�F��h�q��^���wT�a���%�9�n��?~SИſ~�mu�OlIv�4'sT���/a��^��9��*��G�Fh�DM�_��CN�<�_Pg��O5��}s�%��m�o߫R���X�Q?��dK�Z|:�=��yv�k�7`��>y`g�?w����nyh@G��o~>r��F�Ori��)7�9�<���_8)������gѝ;���m��Әܣ{�b�o_;N޼�i�u�Uh��*�޺�#fIuXҮ
u����
#�y#ӻA�XQ�hF��SAC�5�4ky�+����c��$$��co�����кT�a�^�$&�,	�I���g'��cl������S���Qj�0�4o����J�\4Q$�C�6r49�PzєҺ�=����+��iIA���m�[E���*t��P�8P6�� -cZe2��ewv"�.S���x��w�����CU��QS��� *}3���u� 6%��^?|�z�t�z5��Ϲ3.���(N��S� ��l(��sgA�nʟr��>�>�㚋���t=��������������Xpch}0�� ��+V�#Ӟ[��cԈNaH��w�q��Q2S�ٵ4V���2��-��cF����W��ۀ\�����8��2;3�[1{՗��j�A�<�+��sAv��t����Hp(��37I{E���J=䗮�"�c<6��l�����Z#�8�Əg��FM�����4���iu�J��t~�$�kw��E���F_���l��}>��Z?�oW�N�G�SV������aub/���sFp�C=��k�_H��Ĭ�7��f�+8vl�'��G�����U_���
V�sl2|AO����
p�����y��/�9��9p��m⬗��.�|�o%wNk�o�Α���׬�.0�D��^� HK��tx���%�o�ї.�X��gX��1&��e'�r���Sos���5~�) /�E�.+ҝ�_�(6Nk����1�D�2K���XF��o���X���x��>��5�6A�|،׆4�4�"�I�=�쑇��]�(aR9āFؚ����6jk�ͯ�=���~
�b~dF����W������E�[���+���{8�)�жu&�]�I J��r�����yc��T2,ֺ[�/�a?"dh��t��GK�T~��Z��o����7���r�e��x���O�gn�i�G��%�%�O�����r�:�$sf1����O����W��m��<+�)+�ר�_4�b���^�r�A��t�ϫ�kĩǒ�Dn���e����/�v��U��)�ಹ�B�c�P-�VV�,�߈^7�R��I�s��W��?ck�E�>���t�,�ZBrB��{�a�Y͙�tl��I���)X>�hH���)j�]�d�!%����'��S��w>�o�A
�iݪ"a�)�U����*4騻,�4;1��`\C(9gk�M��1|x�ӻ�?e焘.Hx���H�g,��f�b�_#�p�(�m��8R��7K�ٔ�~�Pa:����w��G�=�s�)#��XC�NHM�:�F�w��a�P��8�i`�B�Q=1&�5��c���z��S����B�K��H%x�б�e�	�j��H����t<tF �I>�i�Tx�%�P^��+L+�vs�u�;t̑Y�� �$H�ͣ�uE��E �׽�>^}i�V$�؋+���r�]w�ޛ��R��J��
� �;�x'�)���ܡ���k]�rت��N�;��G����kA3�l����w�OO�Q:v����šf1�jz��V�V�����LN��������j�9]�x��o!��v�J��o��6Yc�$�A�!���-���z_jCXn'��U�G��4j�k�Lʻ�Ӫ�n�
�7٤��	15T�b�a�G��W&�(�1�W���-��7S�>[�LAݸ�Uu��M����ǒ��
Z�( 7{�^��Mx�I���:^�Y��g c��v��+tݙ_���9(����0񠩀���S�Ϲ>mZ$
ש��Y?���.��bk3h�<�(Q�J1�K_#ʩ}{��&[)&�^���^�l��[�kz@�%���׶V�VTĨ@3�M/��~ix��y)�`�.5+�\�0d���0C(Oh�H\�qɌ�oh6���K�(�=X�|;d����_�2�i:�Mz �[�K���q�n�c��-�����k����9�� �3��d�l�rE�(�89������"E��y��M�x�[��z��ᾦ�%!4xE�F����k!�i���b!������g-����|��x��.�M�.�6���y�,��=��S{�|r��5!M,�̠���8��BQ�5��v��I�u���m�C"�DP!��������}�6%$��|�[��`M�n�Y���sٞ4N�av+h�VT㒼;�VT6�>;��|Ի6�a��~�$�(�EoF`�q%!�� ��{M�ܭ�lw�|{Ǆ�"�l(�-��	�13}qh&�ж����G��u��-���⌳[F�t�>�)�pF��|��������t|*�_;�/�˖��Q+t9�z���i���T�F����E��M�4ʓbA,��i��K���Q�R+���q�h��������J {(����|�p�k��w(De]�-�|���<�W�^�Y����J2��U$����G,f67l�)T�y��,�v��W̆W������Jz�����ӆ[���McÞ��w+Au<�	�S�J^bo��7��|�(�&�l��n�3��+�;��Rwgrw�hk�[�@�AK*�����@��w��7;tD?ښP91�XB�6���0��ꓢ��o����Mɢ�h�L0�6���Bʌ�7ʪ*7-r0�j�izE
��GZ.�`ġ%���}~!������ ��h�I��A�G#�c��*!�E1��k��۾>iZ��N�4��J��\��4dA�7]U��r�? �����<��ɮR:�y�=���xw��td�uS� 	):|�7&�5j0��S�
�w�6q5���-g$��_o���t��lJ�������l�Jp�����L��7��>�W��ڄoA�A�I��N֔<��`���_^�J>�����WVa"����c�o�Y����� ��(�ט& ��G�Iv]�����19��8�I/�����0���/v,T<�Q��O��j�ƝɅ	����9�r,���@��VM��!n0��?L�T)��I9F��h�l/�j��T�)ɞp	{ӎ��H=e�����$�?B���bv���b���웊+���.��r꣌�˲�J=ñ0+(��䧄��8Ǯq86�9��R��\ۛcR���~��'9��GH�r�.�	��	H�&F��V6�Aq�3�(S'-�-��àꑢ^�7�{�c���bURW��'��Otf��a������#�mY�hHQqݓ�XH��^ `e��?X ��ٯ�k�����������_9���/�����IB6�)��dq!�d���7��̰gf�⣎���Gף���Q�����
`��J�ւb�^LB�a�?�(S��tx<��~�݇��?��JL�8 ]�ѵZ��ַ��t����j��຤��VT9�)���s� �q4W#���W�C|aB��v�������G��<�~�/k�)Ë �{���=�8'HI���d�2����{Zb�A%1.S�h���8\�S ���l��5����T5_���~�E#�Z�߈r�|׶