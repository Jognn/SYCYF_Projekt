��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&��n?��1ů��> K�-� �&�T�Ek/ֆ�\�놭5�DꢘP���+L+X�4��J��#�0�8���������l��jT��+�(���������6�MC!D�;�m�퓊D@v_p��䙋ⲝ��C_�6�Ռ��#�� ���	RD�4D��畓7���vn�H���0���fX����4 �CS�C`{��;�L����li��� y+����FD�p"��]���y��R��K�({� .؜M�������	^5���ɋ��&���&�@*���
e�� �t+���
_6��O<��7f�M��u���m(MrN����z�jL���@T`��M3��c�uQ�Y���%�dD���,�~^���y@Ga��(����C����	��G�86�S$��ɳT�ز8���:r��/y�[ݦڍ#A�����i�&<nU��<[5)�Z�-Ĭv���0t���d���"_���:�'-��d��*��q����_d�y�N-��~";#��������Y��؆���	6ZJnԷW��έ$Y�K�?�4���L�w�Wmiɶ��Y�?jx#*�i���F�m�E����O6T>]i�_�9;�!(��kH7�OS��_��[-M�((��lO�s�$�g�x7`��ZV�E���F��,9�j	@���]}<�ahb5~ãdl&I^�	v����-�@�@���	��!��d��`j[Q��� r��;f�i�.�m+UH7��/OV��c��������l��i��M��*'��?���G� SK�M��H?�מqT'J,!A�h���'� D��G�T�>��tw�ܻ��l.pRu\7�V-�T�V���CS@�ewf���H�*�cwl�H��ϋ��#�`IY�k����_��U�A#���z\�yz�~�cٽ�bl����S�&+s#�V��%��ӧ'A�N��qT�7a�t��$d��]sH8�G�?����i��i6�ˋKl<�O/���	w�C��:�D��]�l9�ތ�G6���Ccyg9m��<%���o�m:|0�\)!�)�2�*�y�e�M��%����� w�Y�.���,���E�ٗ��N�*��O�zP�i8:³��v�\ݏ*�P�?���`�l��F-U=7�g���w��ȩ��$���"5��!������{Kh��������k�$V,[No�"a�K��H��c&W���Xu3ѳ����i�uI(of���p4<t�Xzf��4p-h��,����<��W%P�)�������c�%w]������"� �ۭ��9�[�Z_���K���N��� �{����Z�@���k}]�s�yR��݋}�k���/���7�&�<�V�0��dG�z}af��5#8��N1�M ��Tl}JĖ�B�	�}E�}�A�	K����D'�R�g��=	������+a������%s,^m�����Ԝ>�m�����?��/ ��#]>؊uN�\���0}�ڇ�T���cj~9�I/g�~0��1���'`p�4��w�:�)�W�M�^�p�r8�^�XO�>j�̫h��BZ�T:�x��z����p<xͿ`����u%�����HM��@\�(��'��b�#d�O��b�i� �SY�L�Z
�=,��H�G�tu�>��^<�Hv��o�z�@�(&\����F��Fq� s�SW�Gv��/������bE���9b�g3D
�'��}d��s�3�KZ�+J��#ӎ���<0}����@A�k%߽����ș39���G�Zx��+�q}l�C�\��xC���#�Y,��7�3��#L�=!¬�#!z6(��Į�bJ<Ρ?�ο�k��kC�����y2<�t�)�.x=\��b㞯�]/�B�w���U.@��CA$��J�0�m����2V�usN�W� �菗S����CC�f�#1H�
�y+,�+��"
.	��������_�R c�Fᪧ�1�&�?E�L[i��4O������{��S���2��Ȑ8��|^�3�]!\rz~n�9.�G�� ���e��	�|�t�?���)ܘ�yz !�"��
��������1W�h��.�R���������,8�Qg�;<d�_�w�n��G�p���]�$�t2����,�<MHi�z�}��ǵ�����w3zT�-Y�%���Ω���ˀʾ�%$���/�W��D���Io��Rb��p�~���yx�Ly���o�$�$?�����8@���
c����n3����|��bπ�����NBg[+��f�u��_ѕ�&m@	�X?�H7�����PC���.�IFc���qs6?�A��|}�_���!�&k�a@o��k��r��3Di�0	J� ���3�6�|�Co��?����)M����|�xƓ޵F���kAضO��@Z�8���t�M�x�MeM/�3
����7�=��R�7���߅�����7���B�)��zݴ�
pN��c�/J�-�G�XO1B��q2ΈS�f�A��Q~#��rӜSY�Ϲ~}g���E0aN#�3��vo�cĿ�'�'�?ݺT�9*��v��_�Ȧwv�A7�oǟ��瘲�偒W^:��,
"W�d�% n�݁�`҅I���e�M�S�	[22d$��ڹ?� �Q�p[���D�fz�8/�qTrĽ$?ۍv����w L͙Hc?�=�w>h@�.�̻��t���MN�'qz&�|���-Άk ��/��hKy� ��ü2�d%Y���4 �"[�g�	���o|;R�]1:ʏ˗�[�������ɔ.O���-�j������[!�[�:"8���hkؑ#Kx��!��(;O�{��g�2Ɨ��C��~��2^c"7��=0��!yc��	��\��=��=Np���-�rx>��۸9V����q:	Vo ��6�3 �d)g'\���鱠 =��d��7�1��%��vBR|�ܜz\�.�ȣo�Uާ��V�9�y�����Ԑ���M))`�4�c%|����a.�A�pG8�FEp��d���e���/�y�l3����Ezs��l9�xҽ�g��IT����ѣ��= I�{+�eP\U�'�]�?_����3g�nF����܊L<���q����X�u��\%v���= �jIV/f%S\e����� ��Fƽ��`���3�o�E�:�4��yc
�	g��2�Jl���6�ې!�*��|3��Հm4eŖ�f�~�#����aĕ?)H�;뜦�hΜ��>�SiwI�y�H��r82������R�p�����
m�8�QU�KkR������]�:漬�NV�����vW�7x�3�>��\��Cz��r�U#_�4/�֚f�̵B�Փ�۰�h��2A ��ҲNR��\�Ɛ��\�g�A�� � ��S�i��`������z5��0�����F/�7<�]�`Nm/3�}�w�)�����hyC�B?3^f��kZi���+֗	f������m�=��2��*"y\���ؑM"Xхu�b����O+�����=�hܱ��;���L�M������ǒȢ�"�y�լ<���+�7x�=��MX�t15��*�?j��!N�o�����7��+ ���zZyuu�^qR��F q@S�6%��T#`6\O�YM�/�����Hq�����:tRR��[^�S ��W��\�MV��M|��e��KX_������̇�޼�\^��Z��DjC���_�!%T��濹���8�����O��mi��*0�"�M죩G'�V)^>�o��g"_��7?�-�V��9>:�쉗��zIڒG�����x��2��e1q�����)h�I@�GAF�]��ȅ	h�Q4���#�3@�۽�j��5H���\��;�ļַ.)�C���{V�W���Ŏ��@�F���y�y}�j�Ax�$���d��L��Sw���ü��l4���<Gԡ(�y�]�9��!H����o��\Vⴼ��G�z�[qC��4�{�1/�k�9H��*�'{�d�a`�Ǌ'~�.II�Q	C����=�z4�1�]_�T��d%.�qDD9{����ki�d�ݚ��w޳x�@5oE�y���)�C����-%����ԹG�����y�"T퍜����� �Tu�