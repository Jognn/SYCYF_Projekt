��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&��n?��1ů��> K�-� �&�T�Ek/ֆ�\�놭5�DꢘP���+L+X�4��J��#�0�8���������l��jT��+�(���������6�MC!D�;�m�퓊D@v_p��䙋ⲝ��C_�6�Ռ��#�� ���	RD�4D��畓7���vn�H���0���fX����4 �CS�C`{��;�L����li��� y+����FD�p"��]���y��R��K�({� .؜M�������	^5���ɋ��&���&�@*���
e�� �t+���
_6��O<��7f�M��u���m(MrN����z�jL���@T`��M3��c�uQ�Y���%�dD���,�~^���y@Ga��(����C����	��G�86�S$��ɳT�ز8���:r��/y�[ݦڍ#A�����i�&<nU��<[5)�Z�-Ĭv���0t���d���"_���:�'-��d��*��q����_d�y�N-��~";#��������Y��؆���	6ZJnԷW��έ$Y�K�?�4���L�w�Wmiɶ��Y�?jx#*�i���F�m�E����O6T>]i�_�9;�!(��kH7�OS��_��[-M�((��lO�s�$�g�x7`��ZV�E���F��,9�j	@���]}<�ahb5~ãdl&I^�	v����-�@�@���	��!��d��`j[Q��� r��;f�i�.�m+UH7��/OV��c��������l��i��M��*'��?���G� SK���mkݛq�K� xwC��f*CU+`�>�zkS}>�����{���K3�&�4�N�����Nؤ	$̂lUPo��t�-ME�U��j�Ì/����$��_s*��
���R�8�Mg7�{T|�{���x�CY�g�"�BO�'YX�{�V���>u*�E&Ҕ����_̯�iz��ڂJ����k���2m��7RH@�u6��$�]�G��=��@:.�D�@��((�c�������X�������:\
��mO��fU��7���CX���R�W����Ȫ��*K	��� Z�������	�6`�4{	��	��#^0�ʄ:��� Q?��qwRK���)��R\fA����&y㈅���}�Kؿȿ[# j�s�N���FEx��~9�?;F�8�6V}Qx�5��dvVy�&E�u2�f)Yk���=D�BvD/r�+ݒ�5�6���N�r�p���nC#?6Aqb�m��`��)��j��r��q���CKr3^ywI�H�S��ڢM¦�-��O����hDf��ҩn�~s��d��`����L��(G��
�}n/h��Ұ�I>��0�%�l����{�x�f���s���Z��v�M2� ���ň��ƽG;��@��P� �f�q��t��L�v���>�˪ְj�A<T���j���hB��'��]5��p�%نQ��jr������\�9�n���{U*`[-I̠@Ix�xm��'d!5�7�֒^찀)Y�4�=(�4��KB~�X�l���^⪈u��عU������?$٫��-W	��n�Q��/���wI:~�}M��{<a} �+:ܿ��ͺ���IxB��>궤
?"���P�!������@eX��]P@k�6�m���͍�L�Ƶ	��f<;�'0:�)�Es�d���t*ưY]~zWad�eXdk���DI�-W��A$��;��h=e����<�
M�^���� "q�3q��%}���ȶ�wN=����Y��v���#P��Q8_gkw�/���Ai}��of�Z�D��~�s�=	P"6R�q��ˠ�L�-��L;	��d�own2*+�;z�a�G4-����8(�c�Ic.��oęy ZV�J��7c�L��T��P���_��!��M�J�݄3�0�p0�����|�kCe�dF��6�C'P�K���4�|���^���������TjX�eSz�;���N4�=�ט������#���|Xn�E�����4�0Pv� v�XQøF�j���o�妧��W2�^^�`���i�)
�P�=���ik1A-�魯��S+�iWK�J��v�Z��N���D�v�֪�(��ve���T���U}�r��DZ^L�i��K�n�b��f8t������R�x/��~�}�\�Ƨ���l.Y$q�ލ��5eY��Wp�Ҷ�[E��`i�Z�$,ޫ��O�Y�v�'aoM�à�N��:S��Qp�a1@↲����l�;�!0����i�������{�l������hۯcS[��OW<\u\��2�a�pr?vZ���y���o�+P@AQ�L�3���0h�X��&��&�����)�$i��I7�u_v���+���-3&m��H0�ê��!G<��wp	U�.O��e��h�7�j���[��k� ���ƞhb,
��\�n��˄m`[E����C ���������d�����,D�u?��ȇ}����+�Fn���0�K�i�.� V��P5��9����o3.���-�M;Y�L�\;tht1s�|ѽ�����D�G�������П��|�������5�%@���֦A�V�f����dZ�`i	UybĄ�b��4�s� .��~�f��^ۧ��UhT�]�����m◟��چ��E,���T�3�m���=���L��_���U��ҥ1�,O�_B���P~�6�+HH_H̗_��P���JTD��ł�gƗ��9��V�:|�VK��C���'4o��C5Y^�O�0���]:\$���A%'A���:� ح�kI�ץ�m���#��R�h��ۏ ��6��q���&u
[=~7�\� `\��ʈ
�u����R�ҢM��X�Z
r |6��]iP�ۉ�d��M��kO�S��iڈ%�~z�FS	�o��O]s�w�a�C�y�5!ԏ���q!~��=^�y�܋d/H;G�"�S�KM4fm���D�K���@��N�R͔�	�3����=:�k>N����mր%�pzD���S�z�v�>v����v�����V5SP]@�Z_i����4qף�~���CgF�3�D�b�y]sA�~��LN�dM����'5� m��gQ�@̦�8�K�eܴ' u�Cm�Zh�b�՚FI��)�<]�3G�`�芷$��f��'��܆�&��6o��ܓW`�����VI���)�٧SZ�G�V�D��.m�_Dk�ɕ"�����[(�ҳ���yy�d�R�����	=����U
��w��e�7����+�tM��-�w�ޤ�+���N��{�_�.��K'�@f᪴��Z�W��|u�F7k{�Cr'RF�0���kG�d�˷ޠ�/�Ed��W-wOA^(֝5 �+�H��q3�-b.��P�rW�����#�%W�m>������7�� ���!.��̀i)5Si�a�q��9В&-�fS��S�^���� �U'WB�H�e5V�i�b�K����z[�ൕuD�r�N����a㖉=m�P*YZ��6�#��ő�Z۽���?�|I�Czhv�؈�?�X@?e{����@E膟̳o|K(���=�	�ִ��pА健2N�R����ݶ�	��W�
�"�o��h����Gm�����=]F�F�?e�<�$l%{ԣ�]"�dW�L��r��Ӑ(���D'���!��ꔃF9ܛ3�
!�-d���[��� ���{h	Y�D�w�\����-�'u�#AH�?b7'�}�1���	��3��)۩ӸA%�%�O�p��.�Xl	�Xk>�q׭ו�g�i���à
L��xf%Q�n���Þ�,nġ���O�K�KÖ���^���mbi���i#��o%�1�]��S0�TҒјQ���Cw�z����//�.��-�#L%+)_
�����|���l�U+�iq>�}��� j?P�K��
2���Ƭ5�+1A�f���*B ��>@�w�0��1�À��+�풛GO�+҄��L�	���{�#��t���:��KuV���=��O]����ul�A.?��p?�TS7�P�x\����i�I�pP(�iuʉ�fwE$
�~��eT�M|2M��D�E���͚�Kkbk�A�ym~��P����a?[;�(^����e���HS]5/Iښ��;;�^V1��*�˓�l���7�����K��H] ���z�����($0Lc2IwOIyҷ��6�z�bCc�0�bs�<�����2~:��FI�xQ����j����; ����aI�����JNE˻��n}l��G�n�דd���!��L�z[�?�:���o��a"�@#�K��Δ��>�tg� 7	_,]�P�B~5H���0�KHkn#�KOw!&>7XG�G��S|�з�#ܢ�'�a��[���n�A_�>+F�d�@ׅ����z	&���dh��t�B�R'�c�h��CN��c+��=[�qS>JQb���}@^����ZgM��s�1	�{�Ml�8��Դ��Y����)�;L{���I d��}C�$����J�ܷ2�P(��>��r�B�V�l������8�'���6WV���:��М"�{¦�U��0�Q<��\�*W|nW���ٙUk����˕��!^4
 0��_JjpV#����*H{eM��0P��Y��u}��,ζJ�,a���R2�]`��mؒ&-7$�,L�;lv� h"��de�f(W�������6Y�]@�
@`�Tc��	��啼�1�8�?��  <-��g��!���d�4�8�1]�a��$b�WO�l���v�L�0��"fpi������[���^�c�F��<e��?����s�Op�N&b%�P�>xo�5������b���Ɇ%D!���z>>����$<[!45��_��	�c��;��N�iG�zrn0�'����4�`�gz~ɐ� �h��Y2�H#�[���S5�Ɔ�����p�ۭp9��S2��rY֌O�>�8(m�_+d�F�h���SAe-�rvW��tdq�O�zL?P<H�l�Da\�:+�ʧy#����Z%���*�$�)/���p��S�aB�N�@T?b��_��7���Θ�
>[+b��պd�b˴��:4X��q��59,d�^��%z"�?���DsB_�����Ds�4hD�#��{VD���U�U�X�M��"��A��A:�Z�>uv�,�)�][���T�<Ą�D�����)
5U�Y�hв˦&C�맫�u�>��ɠ-�?@�� )������*M�bJ�u��?]���¥Y8��)�C��AGdrf�?QAM���\:�R1`q�"g�S��0S��]̨-(ʤgFU!�.��1Nt{Jop�����uu�O%��e}�qн�R�#_�G� 2��0-�p�I����n�L`�>���Y��r$��2��w�:����y��h�(;z���̥�B�JJ�mO�"�g����y�F������!�27�n�ַ}u�Ip��w�"���2�q5�UM|���Ǖ��r����;i�Bɂ?"�ʨíumˋZ��F4�aq�YM��=�Ui�Fhs�PI�i׵�5�^	)Ic��/ ��1��ioQ��{�&�����IXĄQ�T�Cjm��G�xN��'��-��(oAt�w�s���ߴd9{Ƨ���t�=Eli{ °��#d΁��踢��t�`L��q������&�2���������L�e�a�Eb���j.q]� x��>�_�\�(<�:[ ʍ7���f��9K&ݚĎ���6�km�m��`���YhQ����ނ�"=�K��w(^`�PG� H����C�L��?HB�"X:A�zG{M�E�Zb�<.����ĸ�̻�:K�V�<��+�^�����(g�W$�4��x��F��o�U���E�TDc��nD��_.���UW��f}o)��>�4:�W"�Rt?�R�Z�
�|"�%t'�bRޕ )l�uMo�T�M�"�N�����[I\�.Eǘa(I�����7���:�C_�Nm�Y��\����}���^��c�)���磴#V���4���Y�R�m,���윶��Ka'՛������j4�����k�qNj[`�V��Z!��wNZ�� �oˀ�U^z�j��'��"���88��^Dm�%�R�e�%�p�!��-�� rh���q&J�Uð�4��$(l$rh�Wi��	�20���Se��y�M�SrW�^P�:���0�M-[�qZ�]L�jE.oR����}�&Ӭ��M6�a.��H wZݴz3�b8u�����D�%9�0�m��^�����بu�-}�gg��xUh��z[y�d�b���/�Od�IƉ�# ��8��Zd<�J1J��A��	>U�T�ہ��i�a����F��.�$|}L$��!.�Z��=E������	xzp�D�D{a��D��S��z�!�Ƿ�孌�c>"f�L7q� �� �&��&����v�[1ck��7�ˢ㑃��w�[H����g�����Ў�ep���n�>	�j�6�2�[���/L}�9�s����u%n�-2�h"I�Bj��5R7��UV�4�=(^X�T����`������y�t�!K��!��l�޹":��}h7g�a�s� ���I�az�
%���A8��]�����7����|Ժ��e�Y�WG#��я�s=r{ �SOur{O 3�������~w�b%�Y�_do���ۙ5D�=s����BKk����_�u����$�v �J����483��tK3j�'��n{��[/�7�H��z%�/c�L���)<�Fg��8df��[֝N���Kg��@�_T��٦�@���T��E2C�To[t�+{�Ƈ�L��8	#L���X4p�uε�j]Bg�/��Y@<�/�a{���f�y��$����%u�6�&ס�(h�ubqP�4Ca-~����R�W�����g�E�JTA�]�mB�R�c���"�T{��A�b{N���)v�eV!��R�_��?3�*�L�HMVo�[R^��l�!�,J�sA8Pbd�y/��l ���J��|.��;����?�5���@S�
l우`j��S;CGb�T��"�BЛ����]�$��.$���S��gFq�5qQm�\�1u��V�-�i�|du���P>�(����*;'CR��B�3bG4p��-.�l��ϱ�
���;Y
��Z/�{,Z�����m��h����n<ƻ��`4B��H6��"�v_\?�Ƭ@��-�h�>�=3�c��:@(��X��.�*QO���D���n;�@ǖ
Q1�4�|s�>}-O���h���w���'��P����e6N���; �2�λ��M5SҞ���D*�
�����@� ��6�wm���Y�؞�L��=\(!Ύ�9?�_m��n��lz�C�N����a����g8\	�>}h%���b�wvZJ���N��%�kwSI��|��! f2�,׭Z��m����͕�QJ�>�a����0��O ��! ����N� c�C���g*�)I�`q	M�=����Ç��xb̧�@n.������ԛl ��t_n*����` $m�����2����Y�����I�ՕF5��$�c����-!i=d�(�Y#KQFJ��rP���r�΄!�%�
��78�;Oq�ɧ����L4�>O�E����S�NwaJ*�0�O�Nba���xN#׎����X�����CD�
�Ⱦ�HaX�qS�%a6��ؐ|�lr@���,�͂�?2�H��"O>}�7F���>���X����J&:�W��"	P`��¶�tq�Z�͗k���N*�p�]�j8ĆW7���Ύ�bJ��U���K�����m�0}��N�9��!�{���=�6"�1�T�kco�RM���*�X�p��h"��O����Ȧ�{�5�̆���H5��E6�	��'\b��U����g�(C�|��Y��X�c?�N��F*l�����HXn�%�
��8a�k��"15��z���El�1�����-����W�A�ˆ����N��Q�I3'�����C���Y[�!��f���=މ�:��#��V�5�%��Z��ډ�,�Q��E1�u��ڶ�{�{�$�1�*{��n�.��+η᷈����̂D�����[Je#��cťh��J uc���1�|R�!��:0�Qs�*��_Y���|'uL��de�KƖ¹G��@�n��m�eVp�K|��z�(>�	��dfT�U�.1oNj���Nv?t�l�9�ȴ����|h���|���+ ����$�۬��������b��Hz�A�k�͸���z��;�oP�>�.g%��������W}9=��+	a/�5��TX���^�L�#���s��[�Ο |yk̜���D_������?��#^%�r��ƫ֢C��g�����ru�����![ȩd�T.ұܒ=H�q#�4�q�C�2g��l4��P���PA�؀,�e��eA�PA���ѿ�G�4-���쬺;C,�|��-�������n��@�S|��]6�
�S�%���-`��.�A+��.��E3�
��Q��a���Lv�:]ȯ�!�}��}��a�ٻ��	���z��9��s�!T�"�fʦw��-��x��R��~�9>�6L[<@ j�E *�0,�Xl��K.$l��fĊ6-#�D[�P��1j��!�
�H�AF�,ח��摘l x�������}ڞ��Rmx�o͵x\���p������G�|�yN�L9�L�d}1�=� J~CW�\�{�y'�:�	�K.�W$�a����[CT�Q_=�z"2V�ǝ�G�{>�D�N��r'��������� �6��Vڼ� �u�a��p�?�*1^E�vb�W�F]�����vo�OkA.?������<[bQ�����*ɐ*IV�8�x��1����KT�[��п�����F�K��_\5V�
�
R��kk�%[jX��R/����������^;p�`!{; �'���힋�y%�ދ12(�|:#J� ��o��i���k�Y�^ݥ���G�L�s����ԞP��ޮ�CNH���[y��m4��PK�j�i/%d�&��
��G���|�sj2�9"�����e�?�G��<�'�8UȍW���(��E;�P�#��s6OŪ�L>3<��̿����v��d:��2^�F�^h����0w��9�<�I2��t���4[�7Q���F�TB����"C̛5c(� �2v��%�Fm;�`;���Eq�������hb|��R7{5��B��'�+8���*��q���.|e�z�ݏi�p�ù~$X�����[Q_��������s�A~�,M�Y�KK:W�,�˄�.�ݔB�;�Ƴ�U�2����/�w��Oi�>�\u&�t#��6���1�ADf'��Ʃﴣ���G%��U� *匯�]=U�Y��'��K�Ԙ�$V�s�ј� �|kx2�2�dp����Y< �\����B���Uz� �j��'��DWŇ:���|�sO�������?Wn�&�'�!@�MDla5�^M�����s$Vg_fGV2���V7�3od������+�R�=S����E)R�9uG�lp���jo�p�
�.�~�����>1����mk�/��w�Y�������p��G���DM���$"���A��̏?�s�}�&�F��ͤ�w�����,�K��nZ��Id�������9�*lg�|�~D�[�`j,�ǅ?8aB(��"�s=�W�n����\��A��"������ji��������&A����N�1Ɨ��q~�j����`$*�{z���N�d���'[�kU4d�Ւ4���;�Q�~�'/`S�u�/�S}���G�$���U"���9���t-�[@/����E��h+l	b�������"�̅&sVʢXjd*���n�b&ۺ�g�Ixxî7q3d��Jp	�V1���~�cM��\��p[뉅C}88��8}�C#�Ă8�Y�g�!4<�s��ˏ�S�Q)f�K?��v��	�K�1?��j��'b�s3���	n�t)���)(g�\��M�S����}
���oa�P1�};W��m>B7����Qv�g��'�+9]+m�hB�$��k�HWl�JD��ɉ�N���xl_8��	Q�����0��Ee[�o��d?
�*IV!��bu�9HݴG���ŷx���t�QN��`J��}��#�X��H�����Yݿ��ft�;����������b#34�8l{�#��ߪ\۱zy�ȱ����
a�V�)"�Qa�n9&s&R�@����ȋ)�"���0�탃�� !��xM
�AM�?��k�%�V�/��C��7��D�e�B0��*t�s˺�pR����&���9�d���q�"��1�^����ԋ3�� {W���+�����񷭊� ��;�j�VM��f��벶�0�����̀E�w�+d5�����Zkt�g��ݚsK��Qs��?H�I��-}�x4��lFm���`�O�8oƘ!UL;�2�?��8��R�!CuE_����0�8��e�bfX�}�4�������ϣ//���e�N}��'H�d����d�9bh?'h� ���\
'o?}���	�e���j���S�A�����q�A�Æ��v��h�F
<bNX[-�,�����f�����ܯ'�!=� �ј��C�b�U�����N�i�D#��	!�Ŗ�WS��8˅�q":��(�8����A-��п��4�8�{m#��bo\��=:�H���T�U葷M�����]�ʂ�X@�֢�o�'����mW�"��+�@����2�"z$��4Mߒ���{�Y�λ� ��D�lw���w��,��f5�\%�Il9}���9H[�?ɥ�a��%v�������L���k'i�K���92$�nn���*1pI�))�<�=&�9�NZ�M�(��>2��N%��|P��$����me�U���p�Z�F7��Z�{�����ן(�ɦ-���%���++Z�5����[��y&l�_B�Q®���->Ě�
�;�����.,@}3�*�/�#�o��&;��Ho�G(�w"�.Kzg膂��$d�0c*��%�U�T�:E���m�<6%���x^n��OO��PVZ�t�s0o7&R����i���Ā�Xָ�t�7U�+f���:��f�>/C���3��(S1�^{������Osc퍽�R~��٤���8����%���^�"�����9^5�;2�P�9x���㸨�zɄ�|����G8�0�cF�]����f})_x���_�+���烙�Q��W�
��S��&ff�h1�9���%Y�w�宮����X� C��KAA�F�c�&�SE�0���~_�Lko_���m�P�mU岧�ߦ»0�P��ke'�ד�k2��B�A!|AW/�mO$��*e3��5�O�/ť����Ġ����^���z��D�F."����zW�5����e��꠻�H���K���W�?�I@U#�a ZS~v�q2�c�2��d~o���.�wa�2)��IU�:�> �Kʸ�8�<�!�s��'g�e
�	9���h
�Q�W�g�fG>0�������-����* ��8��W(�Lz���u�/#��Q�-�N���%�}�N/����&ʜms���f�6*ݥ�	^�e%�:t�J4��0pŤ��ly?����+ �+��/k��F�7vA}
���]�3#|,����L�щ�RF��Ne^�G��N��f������+dЀ������~�T�W̼J¾���}�D�.�i�H��8��+�ә˘y5�U��G~���=���T.<H����G�&�&�&I�i4��&Y�6G������#�@���kw�_��<$��w$���b#�aGC����&��'t���h�PB�&F��j%��	�k�D��N{m��kաwG�WP��e�Ŵ+]У$���!�	�ҔM�0k�w�R$�o���V�ڽm|Ȫ����3BR/�:e�Y�eZ���3*�0�p�"CС_G���T1~���;�,��2��ʂ+�x�G�ob��p�K�-�SJ��N'�o��Xm�J=d�a�0w�ؠHw]�EK�w/sگ!Z�o��;����9��b+{s�ӆ�ؔnV�����r��;ק8��Qu��Ӄb�
?F5	�wTY�%�X+ތ�i���j��Hq�I�䎦k�L �S��>��V�O
"�����[� L�ޱ|2$y�eD���R�2�~1���P}�=N/w�_�[�3X9��P�]m��p��'�����d��:^ї�$�5u��bfzF��t�^/�eG��Q�_�Gl�ow��j�
{�7O'����TF?�V ��o4��[+�s�������Qܳz'����T��	�	�
׃��k�L�%ޣӓG�[B�_��^v}�B�f�K�*�Y/��
0Fs�89�J"]��
�=�d�)o�'V*��pn"�$K��b�:	�N�F%�;lw��r��2�����8^+�ױ��k�%���Ѡ�o��$gX��t��NZ�gj�D�ÍÚWWz2�=�0��JL�"Of1VQ�X�K)�@:�R������e����Di2�
xx.�ꝆLsL�>�6���y���ז�BWOWb�<���@�j��0�H�1T�l�t�9Y[A���xL;3��&�1��n����[��i�"?w��뤗�����e�斢k'p���@U>!�_p�64	���/���d$!��,����>�^G��4M����gz�+AkEJ�/�w�)$#(a6��v�W