��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&��n?��1ů��> K�-� �&�T�Ek/ֆ�\�놭5�DꢘP���+L+X�4��J��#�0�8���������l��jT��+�(���������6�MC!D�;�m�퓊D@v_p��䙋ⲝ��C_�6�Ռ��#�� ���	RD�4D��畓7���vn�H���0���fX����4 �CS�C`{��;�L����li��� y+����FD�p"��]���y��R��K�({� .؜M�������	^5���ɋ��&���&�@*���
e�� �t+���
_6��O<��7f�M��u���m(MrN����z�jL���@T`��M3��c�uQ�Y���%�dD���,�~^���y@Ga��(����C����	��G�86�S$��ɳT�ز8���:r��/y�[ݦڍ#A�����i�&<nU��<[5)�Z�-Ĭv���0t���d���"_���:�'-��d��*��q����_d�y�N-��~";#��������Y��؆���	6ZJnԷW��έ$Y�K�?�4���L�w�Wmiɶ��Y�?jx#*�i���F�m�E����O6T>]i�_�9;�!(��kH7�OS��_��[-M�((��lO�s�$�g�x7`��ZV�E���F��,9�j	@���]}<�ahb5~ãdl&I^�	v����-�@�@���	��!��d��`j[Q��� r��;f�i�.�m+UH7��/OV��c��������l��i��M��*'��?���G� SK��`����<��M#f�͏H�����������E���5ذ=�bF��<h�U�^/9̰��M`�f�c����\�2=w����'��U	���gL�y	��H���?����,����R���~��7�H��Z��Ѹ>|�,�d�mq��I���%��)��4�^��L<A����y"�}�==YYȤ헻=�.C��߳�鋪��f�ŵ�����#�+��=��搨�JD{<$�*&=�(��ك���E����U��oe�v�X�OMj����.o��~�.h��B�YX_��������wt遵��z�w��vw'�	ꄈLڛ������D���랂��-��7�#��^���c��ɘ�����m��X���e�L�v"��851
�Õ`���r��~nO��k�iU������T�g�������J ��$;�].@{��S&�Gm���۽9
���:sREo��Ts��`����p����iP�N�D q�.�_��&9�3c�
����50�)�[����\N��l��~���WƇ��?�&�� �ST9R
�FG�� ��V�G;�鈤=o�(;zElσ����RDק���}9�}f����N��aĪ�1����}m�=[S���J�/[�X����a��<���� R8_[��ُȩ}�/6�Tֺ.asڷ�s���e��R6쌾L����J75 j�Op�?3�Cy-����j���F#s�Ø���Oؔ�BI��r��P��i�=�j_'���ވՖ� �+�����僚�'�-��*]I֣��mF�`��w�#������b���N-�����rdΆf�E������?	�f���)�