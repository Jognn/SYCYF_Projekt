��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&��n?��1ů��> K�-� �&�T�Ek/ֆ�\�놭5�DꢘP���+L+X�4��J��#�0�8���������l��jT��+�(���������6�MC!D�;�m�퓊D@v_p��䙋ⲝ��C_�6�Ռ��#�� ���	RD�4D��畓7���vn�H���0���fX����4 �CS�C`{��;�L����li��� y+����FD�p"��]���y��R��K�({� .؜M�������	^5���ɋ��&���&�@*���
e�� �t+���
_6��O<��7f�M��u���m(MrN����z�jL���@T`��M3��c�uQ�Y���%�dD���,�~^���y@Ga��(����C����	��G�86�S$��ɳT�ز8���:r��/y�[ݦڍ#A�����i�&<nU��<[5)�Z�-Ĭv���0t���d���"_���:�'-��d��*��q����_d�y�N-��~";#��������Y��؆���	6ZJnԷW��έ$Y�K�?�4���L�w�Wmiɶ��Y�?jx#*�i���F�m�E����O6T>]i�_�9;�!(��kH7�OS��_��[-M�((��lO�s�$�g�x7`��ZV�E���F��,9�j	@���]}<�ahb5~ãdl&I^�	v����-�@�@���	��!��d��`j[Q��� r��;f�i�.�m+UH7��/OV��c��������l��i��M��*'��?���G� SK�M��H?�ç��q;��)��Rȩ�"@���r��Ml>8!�S��L��EgeH]�8��>]GR=&���C��i�Za�z�,�F��h�q��^���wT�a���%�9�n��?~SИſ~�mu�OlIv�4'sT���/a��^��9��*��G�Fh�DM�_��CN�<�_Pg��O5��}s�%��m�o߫R���X�Q?��dK�Z|:�=��y�U�AVD��s���4�&Q��s����F��������Λ�t�z3����~��η�*�,Vz����F�@��W3��2e��́(�r����������d�t�d����\���K�����P0�p�C�G��2�v��í���-�{k	�U�(5�Eo�暈f*+���Bx��
m�Qs�L�pm@�c|��&WfR$RO��o&'��f��QLa��,;�.̰�
L��핋K������
����E�yaeh�tlS�U�{D|�����7'0��<��{cVv�QB��+�D.���;&�>�|$딚�;�V�����[��=w�C��(KK��r��ӧ�E�|��azHuMД��B7��V��e� 	h�L�"�M@ �͆\D���;�G]�_��9�ye@�Mv�"�D�[2�	p�2�
w9p��Aw�_�I��[�Ë2�iC~�����gg�� u�hw{�"۞:�Ҿ�8B�j+�f�b}'���N�#�
�k��*�E ��$��(�؁�0'��v��*�LI��؂8+c��>�?�v��$N���g)���)�gǤ��K�l��R���v��5�ּ颊j���Me��n�BV�n�җ˵d�Pi�m�"s�[�[Qw�,�J�׃0	�����r��1G�7�W�2�F�]���w.&[6�\h����"��*�+E�vQLv��<xh����Akesv2��/�bn���o0�=��ygA�$|��̜-2�P��hMN��4cNԺ�N%r�-�}.�b�X��B�n�UmA��W+� �?\�q�ە������\بA�X��mfa�a�Ƞ�������m'�Į~⫹�f�P����	15W�c�λ�|��҃���j����ƯOAʆX;��ZG;�+`'X��u���3-y[¨���In��C�ji�rpƙ�>T�Rz���k�.q�~��uÕ��*Z#���j^����J���6�SǓP���o�I���&O�����K���[(6O����hb���D��+���'
����[g�����ٲ��B`�w_�(�W�A?������<������� J�"-��r\�4ą��+����ۊN|;�t[|�T�j��ԂuD1�۵��t+��"Ƹ�ؓ���>z���(��֦_?K������$@P-�������n��y>?Y?A^"�Z73e�ԥgLv��J}N7�[b��ȟ=Om4�v�m	�kK3���� g���LK���.2�Q��T q(�X|�ք����I�@����fW}�%+x3Op�����BNp�8�������ºE������UOx0�W�=�H����*�=�=�5��ma���]kH�Y�nm*��@�>�wS3����lg�|bT��"V�|t�@�&��	g*�4�P���n!�o$|��
W*L��=3	���FI�t	V���A.<��1A���k�m�n`ˁ��+1�G?2��C
~��@��8D���kn�h�����w.�o&6$�6�5�KpV�af9��	 �	�T�RDk��.@Z��rjlM�K�9\S?���Ŭ���˶����4�m�V;�͚�1����A��i[�|Q2\G�ʍ�]Q�o���>5s��1d�c�\?���r]c���4&��w.BRꑆ+U�DY>v�d�lX_9�׮���I�Ħ�K$|��io2~ly��o��y^��fL��o{�s�c�^�ɘ�<Ϗ��~]�.�k�!y� ��I���"�xmL�wߩ�>>;��ن�=�=�)*R�Ԥ�<����*�D�h��ɅR0[���[ˮ�'�Wђ��^6��)��� nq��A`T���fC8A��:Z�����^��Ӳ��B�z5i�_�U	�E��1$�Y�<�P-h�(:���oN�Mk�~��pt{�{(E�L	��z�:�H�R��ͮD	!�j(`�Q�6��u͖���A�z���}���?��M���'��p��Hx�*��9�ɉ�&���x��k�[sy�׍���4���0��^m����[a��ڗ.�M��|+P�y��}�.�\�T����_-�:�-�gU㦃G��;%�A�iaⓑE�c�'7��P��c�BZ�IP�?��c�
��I$KY�&��).�V��6��6*���~;e9�x��;���ܢb�5H!t�gC۔"�<��H�u�@��/u�>���XɋAX G�~%�Y�O��ԣ��Y�a~�n�����|�j�k��|ق+P-�ۻ	�@e�C�G#<Ot4I��P��,��}}��
�Q�3��s:��c7��#"O��˾SJ����o`ٯ
ذ�R�w	�8V�9�_����*4X�8s^/g�[m�d���R�HtB���C_P<��'�����1+��o,ń=\�3(M��_c5��;��B g�	R�MM�Z����:K_�ppע�|
���f��m�H�7��\zJ'��>	��,�u�W�ڡ�����B�l"�`,���mr^���`�.��d�<�;�l�w[(�e�1�÷u�G5U��>2N
\A��4�@�P�P�w��0�4~�Z���T��W��p�O�>V,��X!�3��MoJ��J� t$�ӦGo�1e]ll��:�o�x��K\lq���!k�;���w�����@���m�H;i�_a��D0�ZҸ.���`��}�6��4E�Rp|�p�1���C�x����D ���~�G��^�ƅ�_ �7��=_
QE��E�ɘ�2�)-n��H^�$�9���{��bᶏ����R�������g�.��%�О�`|����ˠ�y�v�l�I)<n�y�J~7�}���#��z#G`o1O�+�݇��"#�%[�{'5'�;��#V������-N6_>W�Z���Z"ia���|:8o�̓�jjf�<��ԷJ���A����s��i�󞑇��������`Q��ӗ�䠙_�FE�󈯐JzRي��H�eg{�xAG���t���L���b�_I0�J�[E0�n�A2<�ޜ���,]���M{hz��R��
/�{�5b�@�"���/�; �	xlr��Us����U�F%�������^H7���(�"�Hk)��w��_'#�����]��HT��&�~_2��-����S�k���l9�Etb�BH��m���9j%��78C��Z[�2���*��x�06�i�a�^N-9c ��.Z���[#��Z/�g d�X/���ܿ�j@�+��vV�2u�v^]d�F��R8H�ב��F�e���������]�������s��dv}OZ*��g$@op/�A��@{"�g���v��Vn����f�Y��WA5A�*� ���Ւ'�ǝɨ.*&#�w��t��j�jǘ��x����E����g�=�QEG�%=�+q���?杄#QD ���ݕ������h����+-T��U )��{c�[�u�S���	Φ
�&$۶r�&�1^G]���L�V-�J%J�q�ا(���O���Ь�������V�vi\�_b�V��gR��K����}�H�f��C��&������%S��z�a
ף-�ޜ����f;������AJ�{���Tp��Gr�M��E'�ۃ7���UIFF�a�pF�vg�fGMt����*�ySc��QJ�"�c�8X���.,Џ��o	ϩ�;��6[�Hݬ�/�����%���(co6�=՛�C��̠Y3JUEK�":ʌ��Y�Ns�6�	��t,r�n~�mff�]�@�%�v��D�b~��|ַ-��=�����Q��E����p�VR����n�=�}��'g��5�"��P=��2j�q���tv#O:� ��Y����/1�ƈC���%�i+̑l�+�pA�L$�NBUw���1e�4��s��2eAXn��@��1��n�TjM(A�>��؄�+�T��Z��oVe�J���s�� d�:i�U@�/�C�2�,��8𵠚>K������>^DS0�P.g���|fM<�&䂷�:n���G�>��r"����)x��5�!P�B.�Ue��m�T�]������t`D�ڨ�%/' �/�#���S���j�A���̓���2U�
��S���t�f�}��u�'����v���O���5y{<�'j�s��OU]X3ᒚhg��Rgp�.�b��X�&AZVͼ��}����A�88 ��?�K�M���'���ρy�kXS��d��ޓ��x�g�@1�׈�J�(�K����%�x����B��910�c���/�7�E)ێh%k�Y~�M����2P!qC�*/(k��v5�ڞ4K}>C���j��8`��������D� y ��A��ג�
�f�zw�ǖ�Ǝ���t�U{5�Oz��p��Uv#B!������0�:���S�4�Xw�5Od����]X I���$�Npi�}��&�m*��l�M�y{!�a�Mf,�Q`�����MЗ��[4�+�Ҝ]>e���gS��sH��#9(�(��
.e�:�4>˙��9e�F��5r/�	=Bre(��O��f�de��o�gC�n+^8�����H*�F��$��T��/���Gj��1�
YƇ��&Dv7�3Y|(�9V��}.8+�Q�^�� $U��y�י/ܷ�ڟ9O��밇���l:�pOM�tKE�HC#����Ȅ�-����H����cޱ%�(!���{(9��u�HW{�ɚ�JMlbQ�J�J<B�ݟ W#����Q(Wm��RV�A�l���ȫ�d}P��W�.���T���?Ʃ|����y�1�(��W���Wdd'�����/�����Vє�UڔhOAҿ����+7*|��W�ǙO���[/�6�GcX��S`�v���&y�f�3��d�ȹ/���9�P�*��%�ţpc!�r�l]��S���K�Ѥ�}�
���B��k=*�Ug���	`	�=��wa��̍�(!�ȇKd!�ZH ���vj��b=L���w�~�2{�L����}I�_��V�p��ݤ+v�D�JZX�b��(��� �b�+�j�t�N!��5TR��ԃ���k��F)!���v�T���R ԍ���sO�%3�S�~
�����d*+ה˦��)��h���	ǯ	d_p�����l�����R�0��E� ��eL�+��x���9q��S������V����jU]$`p�Q&�Dv�L�#"ţI�ֵ���)A�|���gY�?{b�x�T7V�����R\���(kb�y��rw�����|K�����w�I5g��-[wH|�N���2�2cƆ�S���=��_�fJ��Kv�a�k���v��>��U=�mJ%ٌ@�$O�x�x��l �{{�ש �Oy��
4�=NJy�-����B�._��Ii�f�����)�ry1JD���dC�ޮ�YR��E=�=��[V�r}�N��m/�C��7��bo����n;����`$�oNna�jY���m/�~���ը��w�vxԠ5�HT���6Hp�K��i��4W0e�`���WCb02�A9O�'���˧��OX}�5>u�R��a_�X��z
�zr=n������ݍv�q�F��/�qS����oxZ �͈1$e-aD�s`"�iC�������[�n9�����MB<!y���Lb��dډr��M���(@\��̩aߵЁ�G��tNt���9��rKO3��+�(�(#���y��y�&3���>Z,H�����G"� �g��N3Oâ��U�t�Y������@��5m%�d���ᫌL�(���V*�bS~{��UyJ�w�2���7��ѭ/&Zߣ[�9��z��ƾ�4�6Z��-wD����6�ˣ���;�3���Lz��kA$3�g�r�?g6M�36�X�T�q|/V�et��Je�)�u}1�� ��v��o>��4�����O�
��P�ϒ�5
�?�c�>:T�rր:�z������Γ���Ȉ�V�t|2���I�'�s��pB�.�k��T���Z~U^���/j�V1���� �L���æq���A����k�{���-���H�fDv�� ���S� ��8r���c*܋��vo� =��p�R�\bgW����������x�D3e�$�Hˊuz�5�a�na՗'�T�}���Z�P���l�FN��`��+���0@M��`"A0Eu"�p��K-wlR�-�W�%�ﮒ�v�^����{8�@����� 	�c�֎���ۇ�+0���j�����,=6��&�E�Ro��\gх�U~,����@���{��p�ß�߱�� �>��땳�5��k��K�py���]n�]x����}�h�� .3�=l��em���%���� ��26�1�³��S2G`�P�^@?%�6!�4U(n�R���XH\�,�]�-���u$��Ѕr����]TclM�
a<Zݧ$�X�'��b���h\�g�í��g�'�!�o��y%/��1U�A�g�Xx�`�LPg���F|�g�-!��Yk1v�OI�����ư6���ٞ6��k�T_,΢�ݭ	��j��K��_߸q�	2(PL ���!'�����f��JՁ�6�q'ζ�_��޸ʸOI�%�(Q!xrϒ�!�1yjp�%�(va��Aw�pa'������㺤a~S�U�:��{%�:�+_~�.�]�	���ȱ��K(e��pM� �6��k%%k��[��Z(1M��������,�i�2׍k�0b���`\���L+�J*in�nr��1�.T<����a���lK�'N|��#/.�d���g�2W��RA
��S?�ܖ�T�q�H��5qȗ*����t_�h%�������g����zC�+b�C�g�� �t|�Y�q�B�r�X;@�p �!��\m��v/�`iu�q�d̩���õ�|�c �T�^�>�M���	�څ(V;U����or=B���R]��;�I�O9�Ο���A+��>g��S�r��|�--;]�3��4�޾��_�1e��nq�o���1hc�E�H�L���TE
����"�~�e<�z�Y����z���Q@��~���.M��0^QS�O}�X��2jgM6��H �g[���(ۣ(�$�r��'Ÿ��v6>A��G��>I-�C��z���~`"4n�g�[���w%�V�W�t�!��66K�.i;^�6���T��/���h�j����>ݜ�Q
9	`h�M�<$4�#�����ps⣨t��p�FSPH�$����1�*)����ʛ��o�MB�)�S�&��o��u%s�OwO�	k���tr��vj�,�ߜ�6��-�JH�uBMXm��Z�f,��ߞ�6B?E:3E�p�i:�
�Ѷ4���8�	�^�^V>����܎�u���kTh�^����T��Z�%A@�X6��ߕ�|�ԛ�iK�Í|1V~��.AJ��	�����P<A��ԭ¸�����N,<��E�k`�Z�@��c���͕21�-�Y� 0�"#�Dee6������"a�lٚ8Z�>�=�gE-0O���FU:E�1�0$�-ǖF��λ��o�>�Wt��@"F%��j�7]࿱z��ǭ���F��"]?%�
�9<�X��l�j(��}7x�u9q��L�����kǧ�b�����&䄺��Þ�k��"��(N���j�%ب�_����ڪ�Ak��~�q�(^~1xOޤ���?�Ƭ�
%�H�iy��`\$�&��J±����I������0t��{�^�/ؓxtO����4�5v�hޥ��������؀
>藉������2�V6qdR�)������M	�Eo�&=�-��rH����@��'��V�kkw�lCy� �n�g�#��\M�j(H�v�K�@@��k��d\2m�)X2�����L�~<y) ������Z@H����^���������S,+4�&��Kn�:$i�OB<�Ĭ
u_U�A�Ł�����c��aN���'	�!��>6gR~���k:7�r`g|HVy��k�!Ml`T�b�:x6V3�TXС�\�~2gD�ZiA���H$�Xq12%EB~�eV��c�<����۶=��B!W����˷�)�-+������M+����xS� 5�ӣ�JGq�V݁<7�^��T��H/�w�k#a2
`��a���f���	P
Qo�YB"����0�`��\�eZ4����`
�Y&�^���	��Wge ͏�]}D#rOF�زu�s&^�hi�������)��sa)�[X� �H�=���������nj���P�Eܔ$!i��$�,_K>{�RG�o���ѷ��AZ���f�Sh������^_u@x��	>t8~u��S�/��^����Ǉ2�3���o���.Yl\�����d�AuH��
B���>@���K�7�8r�AD)�1*�L�zg��T �d���l��AS�̑��"���vjm�r�k�G�U��x�Mq�i�Ȃ��b#d�u���i�@�����T�,�����������B�6ry�t[�sU�pJ�F�p#��śc�� ��	Q'�
�W����lg���b
�p�O��*��}Yf$M "R�ܫ�]4�/�&�-�{Ğ�G������S�kb��I��jr(���V����ECj�#�ҙ\p|q�ql�qG&f�����a�]Ns�d?�ig�=PU	��'�P}Pel^������� 0��0���E>�	�x�Q��
�R�j�ʅke�L�t�u��ƯB.�R�K�P�?g���ǧ>���z�k��S��j��3>����4��~7*��jJ���oa��%��.19����n����?�:����{�Vw,IS �2�Pز��;փ�ӎSК�v�PEЖ_J��Y�ó�-��T"����3��wN��q��͞�wZZ��[W�^���b/����%��.̲�8ݯ��
b�2I$\�s��ğE�r��#��rU�p�pL��74�X44���ۮFwJ����x�k���J��D�*ؔE���\���N('���ʜ(/� ��7-������Վ�ǡ� g5R����Y���FF��k!���tL{�Bv[2�Z�<��J?7�Ţ�w�t��<�RV�U���-k�]���C���$�zUa�^?)_*r��O�. ����+uM�6Q5��]���� ����%��e���tߟd�ș�@Ƞ'z����Rf���<����)�P��������_Ԛ�h��3�%� H�ϰIQ$�	�X)ٶr]W��-���B�K�\�h�8��ӌ�����I�1� ��B�GEd�-��L������]�a-�IX�%E8��z��1��l����\"��x��d��g�����r�9��V�b�8��w�t�r�ɚ���>F���^O碓��-&L�
�I�"�۫�_��a�N~�ۥx����^�h����VGqj8�X���Һ|%dŶM��3�w����,��x%d[��]��K��C�j��C����ۚ%�e܃��Uuv0DY��uhU/W��4�u���ǂ� �E��xK�s�-�=��D �d9����#�=�b=�O�y�g�����|%t���a��W��F��:c�d? /�4�d=����DT�; ��{��Z�κ�?i=�3F��G��k�>��vº�Yn*���O
-)�#�~�{k~� �Հ��A���.�%�]�q�<Ce�2���_���ksɴ5S�:8��\�?V�[��U;y:ZZ�*:a�������d�G�k��h�J4�܍PDR���{�`<��p��3�c�V�/��=�4s:��z��4� >��AW&�wq��K�%�]�����G�����qkŦ�#�^�:&�a��8�S=��PCĚ��c�FGћ� &؅�@ڤ���s���J�씖�-(�T�e>eezYH�ƿ��{V����]p-v���ư�ϕk�y����Ƞ�U/un��5��,nU{����0��=��J���"�c�g�UA�2F�f��5��5�<<;K�YI!�ed�u�]-��MBv�$Xe�f����Dw��������6�&��q��3��͒G+�h��4��G�'�hNr�@z�wO���ĳU�5L�@!gI���Gf<�]�iC��D��U�
?c��y9�a1Ǥk�J��(�*'�Uw;���*O���(�q�b% ��Du�`�]��N�9�W�,KK�&@g����S\�!�����S`U�����@ ��T�u	#_9vA��cO)��{pً'R�֨�����cg�ς`�G2�ջ5?S?stT�Q�x�ɼU��:^yS��j��_�۾)�X����dHDG���q�d����m:q��=����i��2���ퟀQmk�]O��(49