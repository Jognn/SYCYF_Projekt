��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&��n?��1ů��> K�-� �&�T�Ek/ֆ�\�놭5�DꢘP���+L+X�4��J��#�0�8���������l��jT��+�(���������6�MC!D�;�m�퓊D@v_p��䙋ⲝ��C_�6�Ռ��#�� ���	RD�4D��畓7���vn�H���0���fX����4 �CS�C`{��;�L����li��� y+����FD�p"��]���y��R��K�({� .؜M�������	^5���ɋ��&���&�@*���
e�� �t+���
_6��O<��7f�M��u���m(MrN����z�jL���@T`��M3��c�uQ�Y���%�dD���,�~^���y@Ga��(����C����	��G�86�S$��ɳT�ز8���:r��/y�[ݦڍ#A�����i�&<nU��<[5)�Z�-Ĭv���0t���d���"_���:�'-��d��*��q����_d�y�N-��~";#��������Y��؆���	6ZJnԷW��έ$Y�K�?�4���L�w�Wmiɶ��Y�?jx#*�i���F�m�E����O6T>]i�_�9;�!(��kH7�OS��_��[-M�((��lO�s�$�g�x7`��ZV�E���F��,9�j	@���]}<�ahb5~ãdl&I^�	v����-�@�@���	��!��d��`j[Q��� r��;f�i�.�m+UH7��/OV��c��������l��i��M��*'��?���G� SK�M��H?�ç��q;��)��Rȩ�"@���r��Ml>8!�S��L��EgeH]�8��>]GR=&���C��i�Za�z�,�F��h�q��^���wT�a���%�9�n��?~SИſ~�mu�OlIv�4'sT���/a��^��9��*��G�Fh�DM�_��CN�<�_Pg��O5��}s�%��m�o߫R���X�Q?��dK�Z|:�=��y2�}�.�-��'l�{�����@�g��[T_��E�+��6�h�[J��z��o���)~�� j1�6�2>M��y�\���{x����o�W|�!Y@�ͷ9�,�;��L��U����8�J)J�X�o�߰bM�`�gګ�A?�F�)�u{�h�	�zE�Ϲ���h]kA�O4�{�샺!��:���5���~X��[-�B?�B�L�2�t�KNo��7?E���L|u7��c����6aZ��ߺPM�}��Q�6�1�Y'`�/�ɨ�}���!/���t���Ɲ��(έ(��E�4�}2��[=QƯ
[OR={dq�'�W��J��[I��~Bib�dy{�o,������ųT�|aߨ�y��a�?��D�/#�pG3�.��<Uv�^�NMg'ó�F{K]��<b.��3=�,�"�Z_>�y��VI�mM�u1��GN�ـP3j(#	T�6�U��h&����c���F����GL}�z�=����M4�H���&�J5)=�V�_���x��� F��,�x����g�~BF���S������F	8pa���s���ZFQ���d
�aQ�����%FƗ�����������oƋ���5�XrJ�IT�̼�Xz�uTsֳ/�<=*d�q�`�!�Ӿ{-�lC�����w`	6��G�����u,�K�1��Z�aڎ�P5o��-r��s�ǃ������r�6Ut7�* �T6";��eD�-�e�	. 7 �*׹��c�$~�f�BG����oSʤ�u��k/��[LW�k9o���p 3��&kQ9��Q:����4�E���Z��Vj��q�M�l�P�d�*�*�������H��oSt2O� b",�B�]A���b�r�����o|g|�[E?"�p$c�_�wy����s���`��&*��tS;b���jΧ�\����#�?�8�4����f!��7�tX^*5�"2�>Jqd���������oBI�@�6���Ⴒ?���=�0rib��?��QRq_(�_E�Fc����O�UhǞH#X�O��5��0��A(1��M,H�3��y�ss����' ����٢���g��r�����3U��z;%�]���y!Qю�8�6Bz%�{Ib�5�ܡX�.�1}��.$�L��&y5�r�G`/)�?y�^��#������ꕍ �G �F��,��1��L���M��;b�Ȃ���N�9%� ��X>0�ŷ+-l������U�C��*ک�ee*��jO���� 6���.+�Z��5!񎕢�IIi:���Zi�	��it���V�D"��j��bS�P���}�[#yr
g�x�A��N���m�������t��rۤ�ꗠ4%�<�X��{�=M�������P�
��śج\��L{<��=�ol�%�����Q��� k]��ud ������7�S�\�c�a�%?����vj����~1$N�	��\���J�ۊo�M.���8���:mb�JΏ.��6RU$�0��������q�3�f��w�QI���A����:��	@T�2��CN�5��Ѝ��f�{Po����R`�6b�y�^U4K<�1�Uu�J��G���kf�3(2_^������3�
�P��kU)����mKn,�3�q��6A�>L?g���e�������<��I�9�k#�[=|���EN�0��G)Ӽ�i��� ��M��=��Zd$��3t��+�R�2�3h�)W;).	�Mp�L5Hn����1����E4Ȍ������S�0����F�@m 棇n�W�T|�!�Y$7,������,c$%Jz#�
Lb�6�E�.�AZ��J�(x�,��(���$��Ln��TH�g?{\>�:5Y���mϼ��}��� ���M-̓xD�V�Ƀ����H���F�e�P%�5J�h���R?���NY/�v.A*xZ�����Rh*��|��&�7�#+�0T�۸���s3-FΏ�L ���;z`��K��H	��T���!�MH���>41�y�h�gZ�^���5�Nn�r�}� �3`�����`�L� �8��hIuǠ�Qe,�
�x�����ˏ�{���صD�Ttuj0ӡ�*��p$XР��
�  Y���UY�d lR���$�V����-��Y��n
��� ���%/�����&�m�ZoAJlZb�w�W#��ȐM2�x���"aR٦v�4̡`�ځk�S҅�Ix:���&��*�/��i�|�F[��V�YC���n?!wMằ����d�;q�F'��B�g����nN�W��:T�pwo9�C>�{t*醥=P�$��sw+����5�M�6t�RJ��1��2>���H]�ݶ��!y��=�>F����C����>~�#D��#�j� ���u�j�þ�!"^�� x.�j�)4��_�`�܄�I�BQ�ř��I�Iϴԩsd=�&>3-�ay�|����z����7~��DG�:a�͐�8�3
k�����,a~tj�9�����o(黈[E�r��SZ�_{�W�G���._��y���<|�M��?���0Z���"����M ��5���FJ�EB9�h��\{)�@Gվ��/����o��xEb�\c:)��C=xѸ�)Q��4�����/�����).�h��~�)O҆����JUe�^�`�����F�7���i�2�:Ph͐�5�W�y�F�UvU��+Cu����T⸢� 
q�Az����ϒ�f���b���22P�&$5=�n|@%v�t�2e�$0Gu��ݾ�K�zCoMM�Dk �c���%%�X��2�x�~�kc�/��|�xۨ��zZkVk6#Ξ¸w�7����;���t��ݸ�+�ȈY�w��� �5Q 25{�q�`0�?��b������wI�s��3��~	�.�� ��\��]eZv�dq�p^���1��;�I6������=��Nm��^[��b�t8j/�^5ra T6΂�� �9�)��j���>�^ex[Ls�p���؍�+���У��cOK	�������ם�#Ϣ-�����С�Q��fa��%��iQ�c$���a��aX�~�s��VQZ��4��<��#��~�GV�	-�N�.k>������'
�Z*s�Oҡ0��<o ���˛Ϟ
�H!L�Ub��+��R��6bV� (MB��G�j�#rˮ5�H��B�cc��ɡG5P����c���ӑ�+�]m\�/Űs.ې��{4�����<�l�������?��,N�z����y���Ԡ�����W��qJ�v$|��fN�z^�Y}���/X��>�#�-�j�Jv�탮�K�4���a���c[�/E!=P�FdWqb!l�����d�e�<�(%p��U�6K��[�Yf� ��9�֞��Ʋ�V$c��o��V�MiN�<��g3|��|�I��;��Pd-]B���m��	��􋕁�B��-�:��a�b+? �8�F
:	;'�p��)�5o����>���뤪��Hf��^G�� �P��\��?�c�/���H�L!�����e�.ai��2爈�2��u��b
Dg��eYK���c��T�<ۡɧ<��n���P\��P=����:6��uI�⃵X��� Ƥ��Տ�F��H}S��)_���9�|�q�v���}V��2��L�G\�#���Z��n�:�t�^�2���1�&ԃ��m���kpر�"�'��!W8�#wf��I6U�����X� J�v�uw���8�
�������w�9�E���G�,ף����U�:U�̰�0r�9�lc���d{�c5�A�3�{9��x .4	"�:�t��BA�<��ڣ�Z���r>��0����tĮ�*͏���_��b�p_^VV��L�/i��I��b�4s��&be�mv��vm3��Ŝ�D��X=]ev6��	��s���6�K��nC �:ɾ�Σ�/���P���z�5.��m��PP��o�yyԎ>ꋝ��I������/kΓq�c>�o�'Bּ������)�Y�^�^���W�1��I���2>V���n�_Ĺ]:��Z_Y���\G�����Mf�x�b$²���� �"o�F����C�?Ev�%�\�!�� f�4����ع�	i�x6������]o��4x��9���="u�P^��Y���>Ƶy2d5"D�#�y�q�j""�$#���;ĿLpVg�L�Ǖ�$����`X�B�^�A�W!���=S�OM�����%��(�Z�)�mU��V'&R9k{�
�~���`���i�
�P�	�6�5_B-�o�í�^]i��N����T���d1�Q�f��n ���;���,�>�C��'� ��DwOV��S;���'�j��_>p��o׍�${��f��h~Y�Y����ST�AS�$h��!s��|n���w�&b��.S2�h�@g�0�}�9T�f�9ȂR��j�&J(O7[>�y����e��V�l��u�,9"�G�J9�����<��_\�{*
Yc�m�����~E�-x_U5WP~�;[�͂[��6��s�c��!��a/��s���fpQO���|�+[���;�6���G���d̦����/��(��H	#�r�r
�����֐H��c�+	�o�|�A�]��?1��3k$Φ��9{bx9��2�A 0^�0U�?6	�R��Rr�m����̃��]Zѱ$�b�V� b� 4b�{��]+g-��2�� ���O��4i��3Q���J����z���-ğ��v fx����܅�A�-��I{��QH��&�Y�6`~�8E8t ݆�=IN{/@B~� 2w��������w�ud�)ν��!�,�u9�gɗkvK}�<���;N�0����dj�?I���5.�d�*�f��������`Z����F�t���R�(&_j�!��}V�0ktO��JǗeA��~/��"��a�#�k\lD%���͸��[�έgo����tz�P�c"�0��Mg�q�0����]��q�V��𵘎�ފ���ɢ��]���M�VT�R.ڄ��{|� ���;�Ѓ����z��bD�%�]=dL���i����G�7����[��6��0�c�,�(j*�����y�T�4�����\���wh�8]1<�'��^�hv�%"��e�쀝p�ty֦���NN\{e���{�챘M���\�q���K��1s3��'���&?E��ژ|Gy��2��1����9:�0�=p,M�c4�)G`]�O���{p���Ѕ){q_C���D�̔BF�خQ'XC�vns��4�����������"�B��^������Zǽ7��<W]������E�!�}����N���+��_�-RR���9*��> �1;vZFM�`�8r��[���!VMlO\}����}���(M
2���F���Y�m\v�/��Y��<��n���!�$��F΀�0N;ζ�醶���N���X�(8�UFx�5�Gy��f<��D��^i'h8VON�t��^�2�gx�X *�p��7���M4'/44>�	��,a@bd̬<���C?կHښ�~.�ٙ�#�$%�����*�5P���)(���~T �{��$��pP�2նp6J2e���etD@D��hX$��ke�XI���5
I��f���I�x�p3Iv4�.T4؎|��(E���>&�m� ��F^����KԓE�ۯ�E �rPw����f	ga;Y1�_,��e��D�ݖn����{y�%o�rm��^�Q��8S~�߂���:��5�w�3�QK ��}]۫�bs�YŲ��b��'��,x�Q�*Ǥ�>1%D0#d���#-���z�v�Ҵ����r�]ѿ_z5�k�(4֯���8jV�����b���5��m�8�_�c��"�8p�U&`7i}�M��v�Il�:�w��l�;�{�1	"�4xTP^ۍ�r�W�퇇OX���.27��o���!��⚿f�jZ��G�Gn|���P����o��=�Q�#|�G�&�h��#|�>�T:�b�,���fڿÏ\~��G&E�3�<B��_�X| d�����vd�H�N�[њ��ڳ���ų�R�Br���/�D��	�O����@�R�=7��+�ז�c��gi��Б����+=ML�U��f%��>�f0��nua#?j5�
�2��e�]�`�1lFjd��)Y�K��QD T����	s>B"�.{.6�*`$�Ml~�C�ж��x��éK��`��+�&���ς�2@��0Z$z�}�I��t�t���[�>��w���
y�
p�K8D{A�s6իɳ��B�\�>����&	WӉL�׈�IraSn�O��ml2�:���P�]��TX���kSs���1�)�!���tT��ٰ��
-*��v�9��v� ��6�Sm��B/�~��|�7��[-ҩ~�pt�GYΝ��ӫ&�"f!!���^�O�؞�)�mJ�n7�5�K���G�6�ly����Ayf��"L"YX������b��{j%���O�[z��֧NZ���(4	�0XA��61�a���_h�u?�l��$8���+�����F��dC����j�oJ��L_*�t��A
�Z���nۣ��%u�z�,���P�W��R�Cb��{s��P�țc([���7������2VHr��&|���ճNZ�,ѭ�.�,� T̞����S�9b�3�"q.C�RqE�g��~�7���]s�l���X��/�fL��4�$�%�Dl�i�A&��W��Xs�k�?�ү%��a�1e�!e��`_�K>����!��Iݮ�ub�v0���ɶKT	ý��y���H��`��n��c�ı�-�ny?�T�J���Ո88X�N���3�7^���){�w���$�.����r?��ڛN�\�3ǌ�����?k��>GV���ނ�c�W1�n=�1��SaQ����59t6qo�5�|a�+<̖�*�H��QϤ����bj'���9��}����z���2��{�?�W�����PXc<�e�{�x6.1�Di��H�����Nס=��Ì�S�ޫ��&�҂�D�9��>�O��|��҂5��2GJl�0����BI\�^[���9	�)!��Fm?�P�e����s�U�YN�+�$j�>� �u��or�4�>���ݘqVڸ�U����:dw��_Svu����)��dS+=sQ���E��Q��]�;����h�1;�uX�a���؂U�(��W�	��i"X��jE��hkqɽg_�i�'��o���n;�d۔�#��%ꀈ߯��V+�������eL���q{&�Ωo9�d�$.�����:r�E����Y���Ɩ%RN���~_�5Y����&v4�T��4� 4��J��Y{�q%a��"ǿ�xxFx���I����RVՃd�*���:���_��Wd�AuL70|s �im��(τ1���nF��kh+�e���e6L�=>_+���bs��N�?�����t�'�$��ڗİ����0�7�)
�s��hrEٛ�r
�M�Au�&����'e��?���9�7�C�;�&.�W�g��R&���?���lWBm�V"8.Ll���h�������� �+�T�oiF�����1���3 kf�gߊ���F���ߜ�)�
(�&��&��+Az�O��\���"g�iw�0.��޼%���t�|&�u�A�~�����%���g��&�!�T��ژ����Z@;ʿr)���8���S�1���<����]/�q�N�)P�pzl�)�7-�^��B�.��3Y���=�D�c��7]�e�[�o�,��L�|7���;�P���2�N ����Ǝ�|g$R�����
)��>A��gf��1�ZdP.eR��(]?�ܬ�I{�	�|LF	`���si���y�MX�yg�A��9�?�|IZ
ǒz�y���fQ!��T�C���^/�I�m}���;�7+�|*F�|�3�/Va)4��)g\Y�ٺ{��f�y����j�u>[y7��>t����]m�?��(�&L�������~��Z�"��$(+U?��8�����D7��b�H�Qa��hb~"��ٓ��� a���G6�e�!�MFZ���V	�}.�;|�O�Bv�A�ev��8"�>���hil ��g���,@o��s��N��� ���Y|�ΒУW��45,�bنFy$�Y,�������r����||������