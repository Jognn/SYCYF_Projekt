��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&��n?��1ů��> K�-� �&�T�Ek/ֆ�\�놭5�DꢘP���+L+X�4��J��#�0�8���������l��jT��+�(���������6�MC!D�;�m�퓊D@v_p��䙋ⲝ��C_�6�Ռ��#�� ���	RD�4D��畓7���vn�H���0���fX����4 �CS�C`{��;�L����li��� y+����FD�p"��]���y��R��K�({� .؜M�������	^5���ɋ��&���&�@*���
e�� �t+���
_6��O<��7f�M��u���m(MrN����z�jL���@T`��M3��c�uQ�Y���%�dD���,�~^���y@Ga��(����C����	��G�86�S$��ɳT�ز8���:r��/y�[ݦڍ#A�����i�&<nU��<[5)�Z�-Ĭv���0t���d���"_���:�'-��d��*��q����_d�y�N-��~";#��������Y��؆���	6ZJnԷW��έ$Y�K�?�4���L�w�Wmiɶ��Y�?jx#*�i���F�m�E����O6T>]i�_�9;�!(��kH7�OS��_��[-M�((��lO�s�$�g�x7`��ZV�E���F��,9�j	@���]}<�ahb5~ãdl&I^�	v����-�@�@���	��!��d��`j[Q��� r��;f�i�.�m+UH7��/OV��c��������l��i��M��*'��?���G� SK�M��H?�ç��q;��)��Rȩ�"@���r��Ml>8!�S��L��EgeH]�8��>]GR=&���C��i�ZV�顯y��?���-�6D��1f�kwte�Pv���?�N��0�O�{C��=C�T�c�D~7%� 9��!�|�)�r�g�K����vd
�]��I��&��|$PP=x�{�)�Q#�	�b6|���&s�l4��ۋ�'&�u�%��}\�^�U0�B7���}@�hB�< ���}o�M~LM1e����N���u�۰嘓�o篱�:`f.s�c�0�
�t�c�Y��du��V�H#�5�a�ɳ1k��ſ��>�E�Zjb
Jђ��R��y򢺈u�H��/F�sao��TvM/�D�Y7v��T$�^���c'Cj�ֻ5� �8�p���>��t�ɍ��q��X�:���1WL�>���\�-3�̒ -3P�-Q�>r��S�alӆ�;��%��f@��<y�	�汏h:��[��M}ǆKJ;����6�S;B?�P%e9N�� zXڹgE�צt���Q:�m���xh8�:!���=#�fX���`p`�Us�G*��͞�NwɁJՋ?;���B"�}cͬ&��/�u�.������ͼ�|7�������"<f�Xr����#���KK��r�V��-N�bH���oa��P��Bz�q4`.{��.������y�g�v��� ��M	>mA������I���	��u0H�eƣQW$���Ȏ{:�� >G�q�������6*p�8�r]�K^�� um3��b"P:��gl��SXh��_������c�Rz@Z������� ��m~;�(����afF��?6�5�7�ęH�8*�����㊯@:1���5�/�����6=�9��Qds�3��O�'T���oĪ�Sl멭�d�h�l���!�Ʒ�kK:(�\=yk{e��"�$0��t隫��{%�t-Y����󄁣n���o��׫h�'���$�{�/�5������z	�g�HZ�'�~��MSq�gEe�g��E00�S���H�S��)�޲FX���r�F��Vj{l��~Z�6�lA�ն���S�]����� R�f�8�IЎz�����1wzGb������n�|��a��O0@=Se�㨇�(�?<��S����׏�ډ!��}���c	J<
����U����-Y_|��v�cX���C�)ո��@.�����7M��\�^��.Y�)f��l���[ �J+�;D��9�@���-�q�KSS*-=�f�f ��P�@:D�.D�	�q$�a2@��Z�.}9����j�CF��Y�cr!7�!�H��������Ƶ��\5�t�tu���_6I��s#�F��Ar��Fbk��y�G�S)E�$�m0���
�I�}�R��80�#��%���hD�����҄�D���M�H�$�;�z�ʤ�X6�Wa��S�iڕ��С�Wڛ�ș���;4]R\��\.N\G�&�F����-Xl�����q�:ɓ�R!=�����!6A!�;�c��[������������G%:��YT�2h��g���{H��}kq���d�^�Ŭ�b��Ӭ�!����5X�qj�tz�	��F���/ex4;�Ѣ0���$䲮��S$�'��cڛ�����3ݢX��œ4]�V��c�l��&��R��ANe�G��bYp��)�"6�T���F2����;y��"_c�9���;��yKG���ۣ�<��j^eb��A֋�N�V��m`���!*��ƽ �.p�	�Ot�ƭ�ä��D� ��+*Px��P�p��?���"�a$.v��C7�8�v�*��0b��]t���x���X$},�zr2RB>�c&I��,���9 0L����S\f�ͅO����۾p��b���N���Q��W��~���Y:�$�A6ߋ���,e����s�H�P�.z�ב7Q>'�O��}]A�A����i6�dɼ�r5l�P�	�"�WV<�/~��N���w��u�hi��!�B��оxTCJ�b8JP{�p)�!6�v�̈������@o�/H5�y��&qW|y3k:����
]�ؾ���h��������y�A(6���'M"E��C5=�}�j�ͫ/�1��ڳ��;sRwVWJ�\Y�5wb̯�{��U�]&E�cdK���ݲ/���f�%z�݌!}�}#Eř&ZG8�Y*q�s��&F����wA�:O��������L����K"ފ�����E�s�Bj_m��"��HJ+H��q�D5��a�6��/ivK�1��b���H�I]˲�W"B��j�p���գ�#�\�(D�],8c cŎ�%0rD���� ���� �1�:��jo�n��cg������� d�Ae�L�;{��:�"Ce�xV��>�8���w�bqJV��) )�t�楡��V���9Mo,���yC�.�Nɀ�Z4@炯5rK���M&�Pa���(�C������]���vԽ0�(k�G���;�����ت[<�eEW|�T*R>GE�)�I�t�H�S��#(,`7W����� �"�W�0��U��!��Y@|��!|�Y�9rV����S�r�h�ۭX@$g�9�Ai=g�Yw�iۀj`��0��@��I(4�Dʟ���B��L�o�E]Ҵ�)�O��02�[8�i(�G��H�xs\䥯��b@���^�N+Y��>��զ�Zn��a����^�>�P�|݂j�57O�V`:��6fk��$fĆd�`Y���Õ_�WQ�VS�(5X����	$�YY��� ١��&\�^���2��P���38�2����k|���8	ǭy� Y�@�|_x9_m���R@�q�����36��"��|�,��J�I�J����	�g���	G���G��PidxH�I����n�V��pn�_iuY�Y₫����"$z�]���z�u�V��[U��Ӂs����̫ǐ��8ߊ+n�D,����Y/V9`9��,�Nxn\��	7�W��=�?Nj4����+<2��~���"@A/��{0�߿�֔g>�Y����5�1���o	�g�e.�f����c'�&Q�LE�U�����Z��wa_�̱���S�vA��kT�t�<l����0J���:�(&�ƿmfi��0�#�'�n�;٣�3�
���Y�$jq��r�Y���!�>{BB<����~���W[A�4�C�A������~��̶vؗ\�p�ۖ����B�����U�-�w�:?@�-�yd#�� ��"�aA�g�Y�^�M�tt%����t�C��������VH��	��̋�h]\]�X��d/F���ڞ)�����%d�!i%���qz��	�W2�W���+S'~��z������v"�y�L��<�~+�%�������݋�Vl�hX�c����"�1�z..�v�~D�1ٯ���Ξ�é23z�($jZ�l0�<���G^[w �f�wq��up��Y!�*��<�1O�F����U���y,�<��sl'�]�.YCH��8d�!���7���_,o�2�%,����d�H�����<�L���+���#.�P{�Q���d����/B^��?�Ca�(2	��R.�av�|��5Ta��M2���۠��Ef��J��O�q����@�fl��~gg]�\仅:[�yZ[!�5x�]�I �3�"��<	~�nr:��Z绶�@�̽eYG��s�l�U\��� 	R{�Q��}
�_�9'�X�J��2�k���}��U�sd���
�!7�����-ǐ�ƎO���
��V�o4���x>�M�4J�I��:0��xAE����6]3�2{��N�j�049*5�.���<���x�?�B����ZZ������)����>67.Y���Bj��`\�?�k�{�����d�z�́��oN��ܞg�q����qB��v�))+������3�<�k�Ue}꿳�V9��lR�����(]�WL\y�� ��I�<�m�+�J�k=�zs�k�(~�1�����x3|�f���fP��j��*'��*Z�ͣ�D��^��i{�cT�����G n(�߱��~�3Y4\�G�?�P"� ������a]��=�{V�Bͺ#;!CI`u�^�w�#�'���������Wv-%a��x-��V����@Û��z-�|��1TcpE:YI3~W:R���=����Ӊ�)���m���65Zx���+E��L(�$�F��|�m���NP^��bx��?N{���Q�`���P;HY�u��̮I��Z	j!��qHVt(�3a'���b��#�?�]������Y���/�G��=���`�M�%ŶWk�5o�U�ćd1a���M��L$bQ�7�S�,�w��[y�&a�-	[4g�Gؖ&��-\�F�ʬ툌�-�eջ8 ��h> �1D>_ar�Sé�$p��'E���f&����h��&#F��n�D��crRX���K��7��N b)=��>�ąU]�� �8�V<dۓk�~�� ;���gT�W�H�j/M��>�6!�����սL��D�󘜵:���X
��E�9*[��e�}j��j��<7U#&���ߜ���VJ��}l+��ză��OzO�X�e>�"~V\�����w$�X�M�}�H��d�שke;3���e�#���)�VP∮��xv����?&N.f;��87���yf��AR���Q�#>�ԡ�������V�*�7�d�{��^>!�;�ռ���F�}b�qнaB�<�",B���^@�9�y�#��GѴ��m����N�������S�u�T?S�7��s/{뀜S��[����E�N�>7��H��P������[�S=����`2[�]�FkG���6I�)��?	1����Oan�x�'�_�1V�����yWh�p�Y��K%�GZ%J��A�����?�4�Ol�S��R#�V�К�ma����RAXS���⩕ah���[�����a2G_Ѓ���@���\��-���)��ZD�C,�h ?_�Ʊ?t���$*ƀ�N�;��e����E-�YHQ�£Z(K���r�� �q<���>٬<1V:�,�m���E`��|�ST�"H��M0
��f��.�]��˾
��YUtl@:Y���ر����9��Ƭ��aQ �s㒂���R���?�����(<�|�1��c���*�u$�*IW;<o�Cx��&����0�u�k*��fUs�e>$E�MCz�=G2٥n�	#�+i!��@��mm����RPp���2#�$I�����n9:����i&7��wo�����(�&x�lgy��KF�A���EWWg�Ze0��zw�$}�~�Z6֣�V�
�WPvl|�%,t	־X�Yc�O똍�l*��&fP~�v$�-.���@@��i��*����trϽ*ɗ?WM���|��d���� V�}�_8�I2��qk�p�+Ɵ_�:cxD/�E���:$'6N���6��'���g���^�$����!C{\���0��D���P�y�M����)l�˄��L>�0�]M&���;�"1a��#� �w5m�<^To��lY�己��*NmʼN�n��H��:�;S��'~����to����H���� C\6����yk�I�+*�ȩ��Z����1��;/��j����0C2@M�̖{�d�3�����B�z���Ƌ���]�*����{�D��M������y���iF�S]�+^S� 󑧆��0*�~�-5�"��rb�,�b��_2�$�n�MĜ��$�Iї�q��D(=^�7���:�]�T�L���eh�.M���������e*�����jS�Lr7Y���1�5/m/�.�A\��À�d��w�|u9͸�=>�M��T)CЫ'X*���uL�R4��9��C�<_'�����E�8e����ڋ���D��=��h��Y}��qO�ŸT��Es��k]�H)\�ӷB¤�q�2��î`�[��#����X��@��6&0��T0�ԷOM��*9��j}�k�+/$��&����o�sSPV���P��:��J}j�����nMM6-�V�h�(ڡ��s3"j'S�n��"�LY����3�����o� �ic��@���t�.�-�p�-����SVg)y�R�s,٬0��5�m
����ZUN@�U����OcC�g�-#�ee���T?�㓻f��"��_}
j�a�� ���J*�K�A�M��+�J<�l��b��)�V��}����zo�m��dO��=�%��8"��H8�(mz�6k�'e�� �٨h�o�]�P5��߼��_*2�	�ܛ��M\��D/�c̛Xdfo���#���^�/un���u� ��b/������}
R�W\³Oh�����~�c����<ُ�������7�� ӹJ	����`k��<
t�3s%��3��*�u�^�a�	���D�R��>/��yc��&��C7=�K��F�H�������	y��&�yw�(�' T������r���i�ٝm:���A9c�<h"�W!󳐳�|N��m�'�f/������9RN��o>.䈭��0tI�� XY��KU���E��b��u%���r0`M�#�y6�b��+-�]3.�o_V|�]��+�y놜��$�rew���
��97d�o>B��J���UER��@��	�:N��<1�&ۨ��c�H�B�f��_L
1׺�t����z�����ء^�9y�`0Y�a�D:|=h�r�2Zh��ɗxKX�Be�&��Q���;�9�=����xa����@��
�m�	���ʆ�A���#~*����k�Ā�?tkz_�Y-B?9�+9YB�"���LSP@��[���#��h��R;|��@Ǝ��N����
��d��4M��(� ?�÷��jv�Z��1�7v��ڢ���>�\������'��ބ���iN�"���.�P�n�$���`ǭL]C��{�+"��
iҊ�ٖ�����jzy ���o�ج������^֊�����V���WS���{yOQӐ�!+�h$��_b޶A��$Mtl������~*^.���Lq�L�k�W�4Y�,��=q��H娆�Dh�zuh�j����b��3?E!����g5Mpo���ؕ��t���'}u�1��vZw*�2t�7�G��C��Hu\��Om �e4���Z��|W2Fx�i���:Y~���8����?	�[�S�7�~�����4Ѝ�脣���;��MX�� �Q��p(C�^%?��<`��o�G���а��K�P�(k���u�6���8c�k���P���]�pC�x��2�aA�\���tMON1����o�P�a����DX$�Zb�:�l�cq@6�]�ujEќa�=9��憎 \��"��r>�n��>��B�@E��/@˘#���^��E�`���h+ьzӌ>��&����t�,�Q�,m14�p���ަ���͍`���y��9:�z0�Q�y�*hKx2}��*��#M~�!�R�dI:�'hJty!2Ec-�W���"��t�^�B�#��e)�:���y�����p_��P���;ݨ��[_�e��lw���q
r��\�`TlBl�CC�<f �h鮙�k/B�p��a��p�y�O;[MH����b��2����b�첿�����u�Tu���f��r��>�� eg���uK�w�W)Z?�Z���O��q���s�Jn��E0�_���{��R�gm��!ks���O ��F���B0�Z�x�s��]���º���ճy'��*Kgw��U4�<X[�:N, ������E�y��`D>,�S�{?fsn$C�3��1��blvd�VD�R�ύ�M��� 
�_�+/PM��X؂
�c 2ԓ�@����6Ԥ~82݂٧��h���$X�^E��d�eG9�i�	�@b��#�m�ltTQ¡,�;���D��r�<;s$����r��Jǰ������L}a��a�l����q���k��?��7D�@��i2�Q">?0Z���ո�Z0SN
��Da��_͸�A�Z��|�&�t�K��"AQ�T��K��IB�k0��0Z{�$a�i�Ԗ6�=Y�TY]��m��� [�%X�����6o2T~�x�a�$�v�	%�-��QΦ=�F�a��l����.���(�]vZ�ͣ x`'a.�N�^��_�����[5����^,�BKX3،�2�`c7��A�G=���.�Q�Ւm,�\���McWD,Ϧy5��RM%�[�H���C�)�8 �����Ox��Ȳ߲��}#{bˎ�#�5
cEI=U�>l3��R��ݤ���z��x��Ƣ��f}�˳�?��q$����kd���KZ@�Ud7�ua�|�'�J�$?����M� N�0��jM5�S�:������F���Q#�RJ.���|('7a�x	Mt�-��-^/W�Ck�G@"X~U/��}C�3l/x2�ߴ�.h�'\���������4���}�3cw
���k2����3$_y2�u���|�*J��[(@Y�#��O6�'1G�ߗ®Y8��Y80�g�} �|��o��԰��=��XvL�+v����>۬�7��e�	C(OT@��}�4h�bq��iL��$DM�ۺ�X
���F�^a�� j�(����l����hӲ�E��4P�gIn�I�DH�Sf�)��-�L�1��Y�8�4U��usY��s!�����kp�[��aR��bf�C�φ3������"�R�<(۞$V��-:o�h���k,&�,�^��k����2qp瀢y\�[0��=�?�I���.{��8�Zj����Vѿ���].��t/e��;k�����ts�M�Z@B������5�}�GX��J �w5����k�|�g�Zz�孳�ͭ`���|�2��Q[�JD�M�����������=�FNҘ�d��zʗ�:�ha���>�L�bM��w��S�N�
jY��]5��a�-e,q ��ޛv>l��>��Tu����/ڰ��t#�>�D��\�ٸg���-�2�r�B!�WK`�+\��g�2�r�'=��z髏�Z����3V}��q��v� m��K���>ʭ�0Mx�S�5��J\OUv�q�Sc1���-�A�%	?���]��0`<OQ�Nl�(�O�&���?*B;����BcA�,�9�D��;�S�I�-�e�YZ����F�P�|���%wt�J��_�5�u*m
�껄RַX������r�4K�tU�X�W���A�����L��E�cp�c٤�^�J������s��J�~�F�� �D�+���:��& {��z��h[�1�����.��OM�udB��6���~[_�O��n[�8g�=g�q`e����3��/��U�w� 1n��z�[a���&?��ˉh#C�~р���9�1��E*����7GQ�w	��du���wLz_"������FTԸ���e6��<��3L=ٰ�)Y��8����A��;$.vǵ�k{�B�u��05*�v�n��v\CרE,�Q/�t-*����ֽ�Qn�z&ё��l}���������t�cr둡�R�:�m�Wq�M����Z2w]����d���Ԅ2]�q��&(���&Hh��
�q4K�j��#�)�q͛:�B$u��c\T�
�Bϣ'�Y4�w��_�v���>5���x���"��/���g2��TCY
7\���K�����蚴�jGЉCb����C��$�o:ѯ�Ω�X�u�I�Z��iY*j!A�&��bw��72t�i#�Ei�np�����)�V:����D{���u=�Z�1��E�J�"�!��ܦ�=�O���i ڳH/��l�I8*j;�?����Ă;������=��bh�ɜdZ�x?$��� �`�yG��'R��s<�W3��>�ć0��S[[x���"lp�9g=O��w��y�Ǘm����FB��I#��/Ɲ�PJ�)�Y���yy��tԭ�\vp���j��(�0��ۄ�`�:{M�k��H:�^���JY��~4�أ$�W�f���7�)�,jS��e��	�u�������X���^nѳ��q& �_��Ep�Ŭ�� ������P��X��S�[����x�`!�C��%�3����N�'g8H�7���@{���]9�����0����`w.N6��H�tr8�\��7�=�ڜ�ZN��1zU����� �m�Ar�F�_����?ʨ�Ӝ`���n$��r�B��L� �jw?"�% �~Q"��y�OI��z>�I�`������,�d ����F���`�����*�r��	z.z�r.ʉ�Y6���K7����7D~�˴�n�eB ���a���t���#�k^�jw��`h����k�f�C���)�a�=$��	���E�P#c���i@�0m!{�����c߮��}���)�~M�IV���ШB������ �vB�<s.���� ���w/�?��-��Mq���FgL�~!�:�x�^�ю������^F߁�M���{gO;e.���UE�$U������	�a�u���7(��&��b��s��ɬю�0w��&?Br3gt��Ȁ���_Ͽ����T�8S`{0j�j�B��#}Y�q6�}b��r� � ��^[�ޫ����IP�-����A���C
E�|�(��f�!�|����ˢi�Ǹ�b]�W
�6�?���Or�}�D�:5�)=��En��lFӜ�ؙ����� ��z�H�4/������E�dg˲CY	c�r<N�``ľ��,`�}@�B5�{G� ��N?�֖���+��hT�r��\�1گe ���{���$��?�ÖG����J쬖+���v:p��!4F�����$�Q$��z�ʜ���Z!��Y|��l�NL��r��,�=�[��2g��U$�C�%-lr!YWz�9�-n�62[� ,��ܩ��Ma����x�S��c�tys�K�Ϝ�MA�$O��Yͪ1�m��B��[7��x��u��%�;E��mo�>@ϴQ4�ۂ�x�'U��4�=�g�H�@��6_��z����߃k��"�f�G�n0�_��9�*�6*�МF��)��n�f"+���O^`(�Tҩ[S��\1�i��*�@�	"2���Ū��#��+�xu�se�O9"+%�i�~��,����w�C����?��X��l���$��@�����k{R�:� eV�xĈ���t�(��BJH�lP�q�{"��<m�c��¢#x�)]!��L��pt�3SD�@@F�>'@���=g����O�'�.æ��c-%��3l����HT��a�]�rL�v<���ڛ�&��bN�*��S����� �	�ė	��y�B�69@gWx@��U&��Q����1#�v�"�@�C�>��.O8�-h�t]Ƙ��kG5�����eWr��W�4<��7���B~}U�Dl�|ŅF�!Ը�}(ud�@�:�����G�:ő>U�� �q2]��΁;��^��#��P�2�726�~��7��'����0�i�n�a�k�b���8��a��uGW&	WFtF�#ȷ��~�4c�U��P�Mt�	I���������J˻��6������G�7�U��eu������4���7��ރ��k;z��6�0�ّ!2���E����_�ޖ�7���p�{�2��b)�����ӑ5�T\�hT"�o����2�D�`�T�Ih�-u�e9�
63��ŐFvY�O�x�#�q�i��	���E�!�#�KV��%]\�rW��ze���+u�(}���������*�yqi}?p 	��L���b�*����u(�F����?�<�咃Q��4�IA���ᥐ��
	q�;�@�{�������\�-7$U|�5+�|:�.IQz@�;̋������FF>�E��qqD����j� ��t�rO'�\��W�=>O�8/��_�0Z�Ĉ:D;�?��{Ğȴ�κ߄[^�:Q��ߔ��s��b&g��X�ʌK�.���~�Q@vQ����uf���b��d�2�Ob���8
��(���U�f����tW��u�J�%���BHm��V�[���Hi7E�P�A�+%j*=8o_�^��^�aD����Z��N��W�_َ�X�R&&)��� �oY�����"n�Ƨ��+��!�![��K6������&=خ�'�t���E�e�_J�ڇ��� ���� ����H?e:��!�@~��#|�����y���q������%ux�e�E��
΂�.�@'ZO@�-ۛ����O��\[k��&���usk�{�='�X;���^�y�{���]�I�I��x�T�p�`6w	M���k�I<�S�Źބ�O�){SP�Z����co��*���>/���w�v���U�GV��`Γ�K;*���@ �#�t�n�3��D��fO) �p����m��Yq���P��0��&�HY�6��2�P`�y ��5%o��yt5z_��FUuqB��݇�V�a^���d̷�v�3f�x�pxM���t�����m�>F�x���Cݢ6n�|� ���� ��H���P����&���$��E�{�&#}3������7D��ʱp���
���ku�_�m�Fh�@��4���M�V�������N�r������r��Sj*X�>���0�A q�=4��s�${8$���E&S׸ `����dn\�X+~�V�ָX3_�-=��*�l�)j�{��g��|����]Z6Q��n �:���UH����Uw% {+�����i�:ǍG0-�/W:�yzId$�mi����c+"�H�k�7˘�=��uL>i%݀���C����.O�y6���>T�U�ۨ!��"=���M1���������\���S���_B���a��:���H�o�b�n9�7�
����x¥����v>��e��9�*�K<�gt����O�,��	��Xw�#9�{�%5�� E�c��;F��,��otuCp�Qh��mٗ�A���vW}�؞����/t&���nL[gy�g�Q���
Go?��WPEܤ�w"�c�s*��|H��L�nE�t�L������͏J�����R��8�:7��$�����5.���}�RXLl��4"�Š�U�no�	~�����'��m���j�ga���F��eI�)�/h#$��D���+����˟:<���<�Q6�}�R	�-�ga�7KR��ԫ�&���8��-�� �B��Ll�{#[�x;����T�O6�UCX��Ѡk�9���U5������Pl��d�wVRg���5
þ�6}��_9�����2�VF�_�n�����hj��Ƴ�2XI�;K�M5'hWӂg�3ɽ��8a�U�^������/����:p'�$���;�M�=�s�w���F����P!�je�Ke���S�0��6)�ԝ��\h��wM��rN��謀۵�nM�4��TL�{M��l�Q1	�h/�>�#J1�D�,�8��H�����Po�R�Aߍ�bTD4`��b�����]E�tl�!	́�NEj�QX�'1�v>���:�n�:��#1aVv,/��=��[�OS�X�8��Q���̸�Sg���m��0��).�!��;��*�i6��N�b��;Id3i�x.ϟ^�ݤj/w�b�v*^j̰�ZZ���\4΀u�թ A�UK�ٍǯ-��>"�5{S��=������=�_i�)�6 �j�t*$�������^����L�.��H̥ͱ���s|�>�F;w��Sis�Ċ�!��.�WR�p�9B�3pxy�cB~w�bԹ��^��c	��W �,3U��5,7by6I����^��cɬ-��j[�Z�3����q�q1 �  v ���&��4r�d�=�ׁ�s��Y0��Uar݆(%��B#ܬ�ʶ�A
�{����w�SdO Eݪ��硄��J�C�I3+h��1�R4n;�9�TO�PT���-j��2��w��E�W�a*��d2����K ���ao�;G%�uq5Y#<��;�̸I;H��ʦ���<�p6�ND|BR����.<o��箹4dO����K��Q>Z$@'<������mjW�O�G���wy) Ҏ0��PK#��9�I�YB=�+�vA�����Z�r���5XT�4���� �`&�S�҈���-�yn��e��B�>��zt���!Ē���]�z6�O�Θ�S3:�M4���3K����7��շ����5y��I�~� ���U�\՘(�Ub>a���.
w����e*ne:�����=9A�t��Y����4��-�����* /z���q|F��A�q7bm<,����n5�6Wnj9 ;KG r�b���[����J����"]�3�ϝJg�Şx3|S��w`��0(�1�R�y�r��+�����2����2Pks��k����$�3�ƘF�H�b�#$2��z�z���p9!��G�����e��1}��`}�R<U:�۩�\Vڐm.�T�s��*)eP�MΨVi����y �W��o�( ;�>��ٺf�㙢�
��U7�R��[AD�h���l읭Ug��L�iA�!��YL�7#�OX��3�N��i\K:�7�Z�K��=��E9�.>}�	��)�Ştd',L�p�05xn����d(/��0�$�\�RO�M������ϋ�S@�z|״8�c�N��N	���&MYxԏy-�+��	�)�T)e�/3�<�ՆO��B<p���,]^tt��UNG" _�*��L���ݼ�
}^�Z�wSy��+��C\�.�̰��n`�G���R��\EP=m_m���?H���!p��[fA>q���1�*X�Q�ܻ�Iv�q�9֡��˒��p6�Mp�f�y�ɗ�qC_TAh:��OG鱙����{���ܑ%V`��	O�3d����eH?5�)I	�����G��Ex���[�������P�&�H��o<��M-Z��lo�������}:젽i^����d�2f�P2���rC6���*����>Ѩ�ӟ�te	e\������$��9�C�7��h��o7t*��d���[�Zz�?��b�@<���8�Լ��HC/��Dw\!qK�6��eU;d{|	y'%~��@�";�Po��U��y�֊���l���H��+����J������v�x�������u\��k$��y)je6�I��J������]
��zGQ7�؀O���)N�`؂;Ș<kf}���fm����Z��LJ�݂��d��!8�a{�p~H�͈"�2_�� �� D#��vU�O�0K-�ș�X�6�#i700<O,*�C;��Y�Ř�� �`��j��~�"zW�3z.F��\��tu�����3���"���P�`��u����m�$� n�oۀ(]��<R1�Cin�Ra�ە�*$���N$ʂ�2b^;f�9�-��xJ�'mc�3�z$��?'!��?_~j�f�![7J
]k��QtS�|�����������k���WG2�r�(rV�r�'6NW�1��a�Sy���|~7�� X�܆'���`落f�Z<-�N,)H�3� ���!|�SvH���B_;�: �ʸh5~Y��Wh��J�u#�T����@��H��
�}�i	�CG���VGnz���Irx`3�&���Ü���=�����`��=��H�y��2ݤ�m���.��o34=��ÿ~��|NrQ�u��pY���$���Ɨn���}�^ޥ�qŉ,9�h�A��@�T3�����ቑ�Aw�l �c5M�/"���l:�o��3�4�ׁI�Y1΅Z����6�ռ��OZN��[��Ε���r��b��B'h� {�����L��b��3߱I��Z5=ěv0{���j���.�1�;�ǍU��;>�,���I���md�����U�W���M'	Gy�=ˢ�ȕ���{���,��{9`pžE��Ծ���O_"��ɸ�N�TVk�aB���h��",�����GR�\�	ʺr�Z�6��[�@Ï-N�x}���R���W��D��d� ��/I�V9�v�G�
昽����n��-9 ؑ�Y���nق���4�܍ǫ�!�������cI�=2���~V6̰��ncy�˚A.(g����(�����NU�^�khg2����P��jvNX�
�b��ME�o�:��*���$.��,QW����8+;��������lX�u)��0�}y�nj�̻\l�i�	�L?K֏�t�Z9��]l��A���o#�� ڦ�(�/�Ɖ/��ĭw�@�^�g��j����8օ�vU��qe��_%�Dn.� ��_ ��s�j�t�#)v��Ê�J���
��xQ���x��X�a���S8�׾;Z�^ ���+�#z�i��D���s��T�V⇔d��VΩ�˹�u�R"�236�x=�IU��j��ư{�~e�Q�U��q�����<��V� �XT���MڐNܶ�v����ȍ?�T$�:%�ʲH�����30�`'`U��=���Rvh�<Z�ta2�Kb	��mf���L�N���r��|��ɘ:9��O� {���d���ٝքŝn���+�i���{s����zWMq$Z�~Ȳ��W�K�A"C[1������=~�F�G���W�#��Q�Z��^�L��������4��md�A����q��*�n�r<�\D*�b�>��cKY
)&'�3�f��^J����Æ�+N�d����f#W����]6���
'COB�^@SO]�@O-��I�A,������T��G�ڨ"�L�n�r��")���p���JV���y�ok���K9t
J)̟<!(�}�J��4Nc���2�W
�@��Ѧ/���)D�u#� �2I&�[�!'�U9.ɜ�q��R���v��S{4��%sv�/�`A�7?O��ٺ	=�����X�o�I�ZA�*7��y���Ca�O4�4tu��s@m�FB=���&��t���x�8�-I��U�D�	��fBA!����?��z)���T��}`L#!�����AX�����>�W�s����-��0a�>�@����y�=�����bq��%u�M����茋#��J�Q�i�X.5�j��l�ȕ&���9�>�	�K�
��L�mܨ`�mye+雞���3=%9���+3�59�K%��QR95���-��#ۮT�C✭���0��Y���}q�E&���6T	�P����3�n��[���w��5����FN�-�Q�yՙ�Y���D��;�F��䢜�"o򒨳�ڤM��w���x2��e�����p�,	F/!Lu��-�㤐�����֤4�ݞH�T������jao�V���A���*��x֗ ����ݵT~2��ڏj(b>��a�v1GvMi��ޛw�,����5�!�z�D�j���(\��X�-�Q�oyꑘ���.�g{R����؏�w�����T1���͖�X&����¢�t��E]��o}��"+�a:�>ck�f���*��Z������~w κ�Z�tK�' Aở��`���!�!h$F?�0/)n��ʹ��`���k�8����hvY�ʂ��>��\�{`���0����\.?;�:�T߅��*�9��SST���9S���f��+�N��[�w�=�w6fe��Ž�B��~�$�/(4&�r�>�֍�����U�O���XO�2k�8ֶ���0�7�!ϫu嫛���OH�<������bن<���@���U���K��V�����y{�8m��uw1��oOն�tӜ��]�`���)g+u��N���l��VY�JCcuo9t$B�8%��l]@wL�h��������s�%�����;q��������]<��Ϣ��2��\o��iVj<�*Y*I���`���_1��d�V�v�^�`M������X-��Ja���v��緪r1�%�R#�X�;Зqw������ǋY�}��F��ep�P�׈7�
�J++�?��2�b��%�E�@*w�p�v\����~ ��M�#3��(~��H���N��(4�9pv��x(����7�\/��G��j��<ˤT-8�F�]�n}&��͏��H#}�+��}���0�&��JpA��xYƠ�W���]Ra��:����qE�x�Xe�i�o跨�q>��&'3n�,K�*3Bq�ʯ~|�4ab%Mr��O�	d��C�*yh8iI�0�كG7{���_YFg_w��aW�uE,�	߃Ț�Q|�ü���9!�3L��.N�#{9#�l��6P�ХqZ=� P]����x�m�ӬVۺ���R��h��"m�����)ߋ|8�+<:>�딓��Ȧ��z�*��_�V6��]�ݦ��[Ð4�U��O�)d�l2Y��7�@���B��6�I;M�X#�����(��P?�h��Q���1�2�a���ץ!��g\����Btu!��eZ�P$2�i3`S��H	}��r�_~����LѨ�5��?m��G�8$����������u��l���s�\F�Y�0�������Pz5�w�{��y�$�J6SX%�� '/��F�I�cfx v�;~��$Ǆ;�s@�Y^]�:�is�N���mk�=|���^�ٗ�@hVq�aPt��:[_'x,[��0_���畐~l��/ؚ=��"��J��Ê�n"�f��g�a��tWE+�^��N�l��ē����׌\D�*^Vn�=�;�=i�@;�ZDژ��R(�JWd86��:��hMĨ.V�n��l�;Z�{�N��`��6��[��H���@hnK���k�a8���v���_�G>�͂���(���8L?2KAX-�AW	ޗJ4헍~���j������e�;�0�������y�I����`�0����F,j�FVh4v�}SR���-����z���0���3Y��� ���4`��Q}Ow���u���Nt�׍�&��k��GXB��(M`v��[��\�M�c9���Z,w[!�H�1�"�KGBwla��2|y%��D�=	1eR6�>���v	�Jw~���R�0|U,��X��r��a��R�T�G@�H�6�e��������-�z�7�����.y�C늉�KW �5"��16�ۀ��P��@���׆�1Y4b����d�M��z	�'���i���ߖ(�L�ӳ彈����h͔+֣i����-����>�Ֆ�����9i�4;������2�G���Z�/�@�Cj�G9�i�8>Y܍�۪��e؇M�@Z�4��C�G
�U �@�W�Y�Y.ޭ��x��2�	��r��:X5��"u���ezLg�c�UՃM�7nn�I�a�2��晀���J�c�H���TQ$dx�Gah�P\`M���G�E;2��^��f��h����Pޭ�ҽ�#�`E,�nG��nr�D�[��U����������*�yr���ٮ��_<k�_���*�M���-��N��-=�W����&f��6D�.���Z�*{z��h�*�b'��#�x�@ �q��T3`���]g~�	|���V)���iK���½eƤ����|hgw��x��~)�ވ�5���Nf��}��n���?w��{�<.�!y��p}��G�'};�Ʒ^��
I#q��b�?�J���w��ZUi����_e���ɚ�]�)����&��.Q���SG�_�>F�q��W�}�$P�"!N$�g]Ƨa<��[�@3������U�o&��zn�Orb-%닥`n�^[K��jy��9�;Ӟ�����dJ��|�]
�I~��\V����<�EtOMe�Ȋ�s���.�|���]l>yth�6vz��������W�;�y�f��k����r���<�mt�@=���}�䰘��[�1i�ۓ�aPY/eA��b���@�'�;�F����A�$��������j�q��Dq/ē�N_Cn��kq�xz���#m�!g��:�U`m��5�sͬ@-L��c
�l��N3p�1E�s�v2fȫ�숤J4��0;������B�ӄJZe�Wx����-�f��9JO�Z��!@xm+���w�����ZL��A!����ت¸݉#|pE���Y&�fbj{1ئ(�:$2��]wa d��*E���7qi�x�,Ώ�d�!qL��u�SOͦ��d�0A��d!NA��ܻ"�D����wzl�u ��u��XD�'+�_{�u% �����UԢ������qJ ��11w�w�q"�M������z�;7�j^�@{mQ[���~����S�wʟ?1�<'d6�7�lY��;m_5�UaO���L�ujz�ơv�p�#L�eTCe[�:-�;��dN��8��������a~/y��.���V�w��12���FU�@F�9��#���u�}#�j�s������%�*k'�gOď�����MF�q�sx�N�&A���jCA�+�iFR�����:�$���oLU܀�rO�M�����뮠b�}Q��4G���>�J_����zS��S�$�@�O��i��:Z����J�Te�����"����s��盪v�Wlz�Z�0 i�Ot�͑?�:�R�쐭��㊻ŀ�Ġ��nL_Q�|#�0��)e��"��}AK���P��5�3���R�(-l�����d/ �5,����&��G@"]��<��f�+�s�eA���Ge��w_��(ϳ� ���D=�81���V���u�jQ�R6��+2��Fx_)/��tLI�k;�@��;R�.��~�A�5%��Z���7��
K��Z%w@VX%�j�x��յqE��R�Ѓ}��M mޠzw�i���X�	 D����1iH�r2bB`ۗ��EP1�z�������l*������d�;J�p�"AW�5���@Fd�i����<.r�,�M6G��Bފ�l؋0��5ޙ�,�G����	�uXo'�x���g7m+r �͇յ�y��~�vG< գ����Y�	����F�D��!�PM����|c�$n����Nغ����Ĝo�9���5��$s,h�LoV������ޛ�O6�صѤ�Qi(�V&@b�t�3 �o�4��b�BΞ	kI�1����0��@���}:�F�����Ww�)k��0��r>�}���u���n��O����~y�xL"y��Ɓ��_K^t �n��,B�s�WR���Ӫ��Av���ϩ�{�+���^TDxb����@9���Br���H�����
`����,2�k%�g�(n�x�6��$(��H���u8�9��]���|���wd7�^Β_�2)C�e��9CK�ž�T������],w-�R�0a�dq��$�m1�2�e���T�˪݌�\��+�\>�*wwR���ƻЙE-4�.�G�5P!v7��-v��X�W��1����	�h��b�b謸��B���{�����+���g<�*�t��&�d2lh("����	�Q�J��|��%}�P��[�1�f;�҆Q�܋���	�X@���~��!a��ݤ�ځ�?:�2~��[s���3dV�^�������LQ�{PO�u^��h���4xx�X��.�?���v���>,~�2+M�׈�K���0�*�c�X~�S���?�ֵv�ׁ��KP�٬][�9���=�o���97��s
��4�%?�~)ے���`.��@k�f�A���"������T�N�����6�=t�+`���g���vqkmQ���*�5K OB�2��F>_:=�4���K]]���� �kŭ�?Y6��2|5�Qo��!��lp����f���%����#�2����\n�F+�/��qx�:턥�ZH���I������v&7�.W�P3z�c!D��A6u|�Dw�&_�3y$�d��/WTN�J��Tk
�������^Нb�RXH:��^���7��x��k�����@�HA�h��P�BH�D�n�D��^������]�?T�  �����p8j�]�3����0.3).3�p��qH�|�b:Wc���N:��Ai�S�:���Q��H���ij��.�0*�0�!G$���x	���6��D	�dGꋩ�jT����-E�U�aC>��x��Ty5P��L�4�x���vv��e�\;I�(�B\)Wu�Z���`�wT���K6�_�Ų�g8�+lH��L���*�p��X�q�(�z�):WmXIt�>')$PC��+�t��\V��7o<<�~Zۆ��bN���%�����T��uȆWCC��_��A��4��M������G��R�gW�C���XK1&�/,��Pa�8��Z*d��ބ�CY����,��c�`�[_.k��|���E�
�Q�iq��)�/��k�;�ب@|�DO�{�!��03௹���؆��o�H�^F]#���uȋ��n��qZo_�.o~�d���:/��TW\�}���ؑ0���`�9��!3�\Vr'��k$[�#���"� �ʝ�H��|��*�g����`���x�Ƀd���n���z�|v��J��P3G��̲�[?���7Y=c�?v��M���/8�ȼ ƽN���|���5p>��N��# �s��Xؚz-�Y\�-���ܶ�2i�E�ҾlRc��/�b�L���I�J��?���T���w`8qH|F�F�2�/"�����_ŋQQK���+�D�T;@��;"�ߛ~d�"�'{�V��1co�>;����\���$DG>̀��W�f��L��mOw� ��yάy4n|'��� c��8P�����	[��?t�%�؎A��]�������QZj��*Ё&�N�&��K��(&|qϋ'E�ye�0����sh����_���G��u����r��E�/�b�wk���<I����x��I|o���	�=z�K�!��޲��l� 4Oz	��ZX�zh��.�k��Ī�:���b҉h# Fف�Yc��	^P�*
b���AW)-�P�#`M{s���ah���n���a�T����Hֻ�]6�W�����iPu�v��0��1�#�7�%Һ�8^���dy���N�|bʉ�1���\e�h��k9+���ۃ��EYNsٮe�ty��ĉ+�cwx��'�İ�,�GV���a��B�O���a�����]�!�r�@�%�u	uU�e.L\E	L̆�ت�?����-`��%�&J2�9�Ԟɑ��|������wŖ�i��F����*�H|k6?	�W@�x����V.��<��"@~u�8��D����+t�2SvCf�'�7R�V)33�B3o!H��ơ�b�D~a�F:or ������c����I��r�l_σ&��Okjv�ɗ��6�ߚ��j�u�]����(��%5�̒�[�$Y������q��!U�����[�<���]x�B�}ǌh~�BQ��Cn���N��A��L߂��;h �z6qt�0�hP���|I׎��6��$+"�U0������o�\�K<��5�)&�`�� ���\�X8|��� �TG�'��N3�]
+�!Yn�=�sc_Q���4+��5A�+F>�_���l�#�;�yX�ޙ�E���=�G[rsH
8���Ⱦ�~Qm9?�۝A!U�	B��!�_8J�x	�������K�1`sPc�²Uj��ak��暵��|�i{Ո}>�׉*<8��,��	�8V,�rdpv��#X�L�t��Hf���/� Q��ƽ$>��Y��� ������eЀ��)�
�H���zڙ���n��E�]�����B/U��1�.Y	+����Z�����(���[�7�.L���\^ k�+��2zTC!�V���#�3��ڝS	������>Gj~���F�R:w���E�d�i�p�wԮ�6^�����S�	����j<�h�*S�xyP;o�h��i(��s�dE���4��}�����o;p�| �K0���]��]������Xg�V�׼��螋��*�dgl"��9w�M����kM@~����9�^[ɵ�gVl^ɤ +�AM~�ۉ����j����~&�ut��f���)qZ�����S�����m؈�ùPn����+��I�S��Eg��/^�
#(�3����(^�7�ZAr[�w��^d:����b #�l�XHJ�に�?��ߜU�͈�!��N}�Am��TB�,E�t��l�%�.0�nH�S|(C$r�Um�ŸC3�(�������@��LՕKA�#�܇�_�^��w�B7��P_e���9ɟ��=��j�do8����2=��;��(X�	��� ��� W`����*=���?3P����ᅂ�E�!��3Pt,��n���+�������(0!���g��E孬��[e����/�7ȸc���fHt������0Se�9PC��h�h���W�e��#�*�/��81c�,>`��i��W\����w�hoZc���`B��n�9f�ط��4N��0��?a�Z���t�-{�E�2�,l���x��V
:��"L�{��ˊ��z���ͤ&��k\��Vڂ6TdoI4�ib��B��������bW�8g)`(Q}����0�Ϩ�{�|�=�Y�H����¢�f߻$���",Htcl�"�7��_g]8���ޢCo����NE�sa�e�CR^��u�@��Q16���ˆ����7W����Eat(����!a?�(�g�G	��p��,V%�b>��8-v	�\�裗���o�HQ_�P������W�O
�1b�������e��*^�Sɨb��C�j�k��@M�p��u�`y�y�%�o�5��\���C!�s�0d^/�����~�J����HO�ý�M߅`�;��h�ٝl��79A_y��Z3ƪ�4dtC�V 8&����A��S��O,ʠ��F�>Lr�YP�����m�XFvʻ �y@��iD(��-�<���T�����,�Tމ�-]X��Wη�_w�l�5�
\����2�3�p��8��,K�A������J3v$2(b=�3�G��p�?�����o�M_�Q���s�m}��T-������S��{����Ƣ��4�|mO�M���D�bl�*ǌ�ݦ��G���=�sS��LZCCj�bqeB�Bo�"�8O)��6F�
I?������#>��5��p����8�"7��?=P}ڮT�6��Ξ�T�:N�Q�ũ"�El��j wmŉ���(���y������r�p�_��n����Kj��C5��=���Ϥ`��`�f�J\��ڡ�V���x8ۿ~T:�"	�2�IM�����X�����Ӎ����
� G�#ߔ��g���_�����y��H����'ڴH�W1	�f7΃Nr��fo'����� ����Ig���YP�.<����r�#^ �/��W���֗@���js�«���g�Do������N!e�m�G���3B�舮V�kKk�"X��/���5Ix=,�.㿁 D����f��(�]N1.\�i���{�B�\�%O�a���/a��>$�t�7����~�M؛r�t���Zr�jȅ=mA����t����鴯��ժ�e
./N\���C�o`Z�H�{�:�<�V��| N]���U,�sQ\vB6��>����	��+!�G�O��!9��>�yXз�痙��C8��c�)��2Z�x�8Z�qW�h���H�wP��j[������t��bw�P_�w����G.}X=���uq�ېS��˖��^�� �b.S�]!ዒ�ka�)��׿bԧ8d5���N��I�_T��>ސ������-ڒ��� v�cz2��N�W�I�B��Ԡ� +����-�>��#f�.���)chs~?�o���a�I�'��T�,��M5>�7ѭ$Bz���Y<:b�
+���J����6U���˷;�M��:`�Z�_�f,^�V#d���
�8^6�8F�����l��F��6=�o�����
8Sr��$}ȉe�1�S���}=��-'����՟mp�V(4��B��᳡�&�D!��{��\�IF��/���UZ~}���m��l�>(|:>�+%��� @�֕|��ra�=���5;}���T�Jc��ᡓ X�/9)��A�K��7�����r-�l��/��<w�QFXe���0��W�+]kx5�^��n5�g�,e��`�}�X:H�}4V �/�6Cg#�j�uDxy@�|92t�C�	�A,���� �c��iC��8�0kI��WS��j�?͛�L��ge�~����&�t�:pˤ�	����ҕ�f|�%���eK�mb(�p�x��Z}�'��e�i�<)��;ڔ�G ���� \w�?#��d��]�Z �_\�OB}���S��}�`թ��kA��h�rB�u&���2ڡk$��A��W��V:r&]K[����(�m<�i ¸����7����,y�$팡v#�� e6�PR�{��Jfb���ֻ���J���X�+(��j���92�_���F#��g����˳h� G҄�\Ѽ���+�kg����d�.'�
2�.��r�ن��`Wƺ����7Y����ދX��p�`h���a�����c�Ѣ�����iL�)�I������e���Շ��JG���jD���:�`��\"���&��cg`�񝽕��
�H���;��V�e�L��Ym����1ľ�u��
�n�F��y9����41E��C���q��)�-�4�O�&�xe�`9d3�14uVs�E�Aӫڱ���"�̻skV��J�Ş}t;��u7��o9�w�Xd)�"�v�P�b͌�^H¬����@*�|�rRL�B�^��?��¨y${ċ;��)��3nBI�&��}��_�Z~݈�Kt9Y¾6��{V<���*y��|CR%�k#Ѿ���`{�8�J������ũ�d��1��U�����q�]wSP��'S�۽�o���TA��A�ٍ�|D�?4�Ud�>�2	FF�=�_���E�ʲT�f��xԜR�Λ�5�\���_!��n�*-[;jE��س�x>��_�KԫB&%S�I S���e&U�V���O|�������b��;���,rϮ�v.�aa�n�WM�v�/��ǰ�5Kg,���O+�`V�>�1:gn���͓?��i��l�,2��1��׶`0Z�P�,��}O�ꉍuG���Fϓ�z\#һ�>�݀HиK���x���c���dU��N\�T
���G"� )�w[t�3d�.�%�Tr��L��
�N�*W�2֞2(�al�/�4?84���sf&�K�����Z#��*c� �Q��F�#��U��fwlI����x!�ٺi�$C<�_R\�[�Ր�,p��oBG5Ѥⴘ>8��Y�/u�F�q��Q-$q�������?���J��J��%_5�#�PN��%�T�̐J�DrP���ޒ���զH��n�~r���]o����#�5=�eI�����zyF|x��0�
>|4����yj�����~���Ep\��[���QQ��U2Nv�[�%���d�I-�c[e"�Z�&Q�7�r<��� ��O5��o��IWpGA�����Vh�����F�8�$�D�F{R}Ǵ��jL(Z�&m�Ou]�ϗ8zS�R|���}���@�I��$w(�B`�d�@Vz��lp���@կ-ʗ]p�@�.��l����ce}V:�t�����9���-ޔ�n!֕�M���P7�O��B�V9Ka�)�,O/G���X���#Tf��iS4�D�y��V6��Rv�MO��N ��k��
3O$������Ah&�,W޶v�vp�v>�.����<��Zo�����S��堓N���������n��OKO�MS��K��xt�v�'[��6��v����e�B�}�,��fDw˺x���W�?$"�[�=�ˏ�5��6o8\�� ;<�E���N�|qX��9J�Ǻ�H��z�M�EC��R��\��;��Geߦs܀)��FI�9��5��YGy�������5���MUB��Z[�"F�!ݠq����i�o��a�m���JPrrf�fU#W+˙�M00���{��V��4o�~�H'�QAB_+�&� Բ񃷩
#&����)|R�� ��~�mZ��P�K���@o����QdF���G�{�WU��_{5$�{ǞT���>��,�T��Lz����B�b���L�w_�ǈ`�v�A�+��J��n��c]&��́�H(}UA6c��[#�B]�&"��^��q�`T
{|6�b��"�l d���ԏųùW��/�8�#�7Z����ȤPpD�>���nx��4�e18�>�|��6�`*���nU=�4�t�47�r�����*Q�]��+S�2S�`V�x"2c�:��A|� �N� ծ�n��.K7���p�՝c�
��RZ�D&��t�v�%�2L$K��\�� ʺ���E���6�[��qx�y*��z ���� � �C\�#ߔ��Q��KiC�TC�/�aBU����5iee@�=j���G	����K.�l!3آozr�]���g�uc:˞3�D����(Տ�q�Y6�\Z�(����uom�S?��V�~[���;>b�1]��bWE��%���$�e\��H,�F#��G�R^�鸩�`�(x�d��R�}AV���	�#� �5Z�������%NY�
2�ф�󁡃|�}w��j��YGR�b����O�C]��{E��͒ˋ�~(���)VW5�L�C�Q���w�_�u0�E��p\��X�:�>&+I�����>�E�9�+~�����UҰ��b��7��W&+a��r�X�����4���ҫ�¿������u d��*��kgl\A�ο�9�A�n$ra�yL�%1ؑ����ݝ<7wΖ�~�`��@�"Eg�����}����+$�fYH~�u�J����`���b�,�w��g�����0�gXi���e˂�v����#����h��vUR��W�r��?��J��p�D<�:����������~��s���	4z._�.��e���c�ERys�`W�Z�-��%~�f���{��e c��ꑲc��^���M�� Z\�4�/kKf G�6�ֽ)�>� �e�C�CB���.dN�6}O!�|�.MJA���:޼��Hmt+3�X�u,�ז^��鼢����/�A�i�[����:G�5�����3,�o���z��#��H��S;������'���՗���yT�׾gu�z������;��Xi}�}��V�r��@%|Q�{�+��uR��9����9}���q�edA�c�����D�90�	��w5P����a݆(�=J@LG���b�@�TV;��������ē3�5�	_�體�|.0�z�lq��^�Ot���B9�w���59P��@���GO�K�<�._��k�m�5䲄w�h�Xs��X�n��	PvF��u{�ߕ�<�F���-%H<k��9t~�J�&K�/�t�Z�s�M�:\'1k���(�ld���8V�|q����w�l��e !P�@Zy0��'�tыE�C�ezw�*NY�>0��.r�Ψ����c���H`ڄ2���ɍ��	n�"xl/-�n�v,-)QT�� ��r(t�k!S�]5�[p�!��$��C0{�Y$����2^�4Vtn ���ʪ��V�*������G<RN{��5�W���E����yU���\�������B.������������[��Rg!v}���֫�@>��u�$9��Uu�ài�J�1��j�Q������T�/D>�!`=�/dȟ���ޫ�7>�)��hݝC�ˊe��#�k]	vM*��㸊7�m��q��V�X��1ӏ����ML��q���^Z��#��ǳ�p��S���E��yz��ڼ#!�ObL[�aV{j`?����z﫩��l��%x�������<u��]N����p��H"Z���YW	0�z��	N����Pƀ��U̔�/ ܢΓ)�Q5i�/f��]aT^�u`Z�f��a`IѢŸ�R"�7�g�{XٮKc-Z�`�=�<aH���V ���w*���qN���,��j�"�).�p��6����S�I�^��'�J��c{Qӫ~�·�:
a�d�l,a���"�=�|�~��q�pwaFH�PĺW��˖e�-�8��J���ns����Z���w�P�}`p�C�ڼ�~Y�=8$uw!�)'<a����6T��9d%U��N#���C��9s�f����3��3�`���tHH`yC���\�,�0H��b�y���`�@|K�`w�op�N���t_K��7m�U߉+�pS��8W,.t1  L d$u�L�>��"�J�;f�'U�>D��Z�B���4�!����2C1���v-�>�}y+�p|A�`�A����������1��`q!�?�*� C���j���9f���vaWy��J���0��WQB��l����ybA�夵ԓ�xơ�X��+$�����RҤ|��h��o���a0Ld1���C'�-����K���?t�=P�Fۉa�5Bը�VQ[�IX�Zd��3�h��z6��k�]W��h�V�2�g/���U6�č�O%����:��A?�3�7���*r��b!`�uR�#���4u!�~�}<>5��U����n�\�E��п�J$�n��X�um+�)��E��X�zA�G4|2�.�|u2l�%r���R{��~�Q|��w��c���B�izNb�����+��VG)�l8�1�r�݊����7�UC��*5,B�Y��T9���hӋױ����O��(�Z�\�o�G��a�y�*���u��|n���?�QV.�k��(�8f���Q��� �����lֈ�b��*yn�HJ�ߴj|��ǋP(\�?�9�����>�B$l6���D��֠�&�N*;�/�J��p"nQ�.���,WcJ�OdK��\B�h�6V̓�/�E!�JȋU�VT��L���k����p�֝��x��~����z�j���뇠2_����Dp����(� �8}�A�?�n�`<'���
\�f�}�u�N��t��`z�%�"�rGl
$K1���K	�Vhq疶x���&c�Y~��3E���Sj.�Y߭����0��߷���=�]9+������mG�1ݏSC��.��Zu�30�Y5�5�8?�|XAE��t��X�mƃo*T}�H�:��_=%0a�M��*��u�����#��;D�eE�1��ٟ�w��]{�DrKF�{:�l�s>�cޏ�Js� ��%�J���(�����g�
�
���x���;��ON+�>Z��%;�"i�e2��B�������ѐ`~S�r��.��v<�.A�T��ߝr&�/!	��/�%}�ZX���4TL6����ɋ�g'c=�5�,B�)!�S԰����ڙ����s���q�+�� Y�В�{��*���h���1��e��8�����S�{�Md����1�-K̡uG��q�v�%e�]֝�i��#u�{oD|��� _��0�o��U}CGS�Uf䒯z���#�=�Z]��-�+�({z�ΘKژ��*�_u-�蟖��ji��!\�g��@Tk���+�������~�þ�~��9��L�Hu=ST���8��5�V,6�Bp�g��h���@:�^�	���	��Cm�!�����sqM_�@o��H�ǚ�5���Y&�R�!�I�X6"nA��s�᭏Q��)���h������ƒ�j�ȑ������J�5�K�y%��b3a�+@v��=��]�d>H�"�]��|!�ǋ����ߦ�&!�;t�|#y*��%��c��|�+��^�6]��+I���y�:����N��*�	�~cҌ�@oqF��������J��a��p���ۗ�H����N�q��[̲������K$��	B'Ȕ����-�~��ס�P[�X��fY�Z�'��U3�saj�3��X�&;�<�� �[�2sJ��D��ag��d��)M��"��q�5�C�gB0+%�&O�=����}SQ��y¹��F�s�Ԙ����E�����OZӊ��7�N��P���6��a��a�&��a�w�x@�3����R\��_���Vb}b�5�3�['�{�G�K2WX'�G�%.����5Oz�q̻�+�.�%��6吅�6ey��)1��K��HP"0'�R��]^dk���9L ��o�{\I^������+)��=���0���݂��V������^���B��,saj�^I���
�F�O�c��=0��_�]9T��֎U�~�����ʎEc.r��-�_�}+�Ne�`�<��*V4G�x����W�����,ѽ�c��GV��v"Uq&��Q��"�`L~v�(䯁D��D��يIg��W�6���$v kŖ1.�(:Ǘ!�6'$�)���/(���r';/�D���-m�Ѽ�/g
�>ՙ��.7n���!��f���tp���K��7�tA8�@��c�j�1���p?�=�_�ɭ�wt��m��a4d{�u���o��f,.j���؆:BI��̆֔*�te5)��{���Z8���m6�X5���5�D�d��'(i�*���Z/���鹾�3�����~ݱ�N�H����Gތ�e(��<�Fh�H��+�й���ɹ�S����S�������W2������&���x�B{�I/�X^L� �v�����b;;;��u1��YI5��	����>X_(;�u�%�	�,�:I�C?��ݛ�ё�{�B�K�eٮf^�"j����Q�1
ǄE��<����.d���\�э����۝4Ĕ 7ڀS]��A�xvB�"v�6�J+��<���|�.&bo�v0�w7�a�l�
�p��1�q�D�f�x�#��2���N/Ϲ�iQ�h�/�t
�ǹ��P8�,��ދx�4�H�9�J� ��Hցx���%���(��ͥ"���D��̋�#�0�~��U����m��Pߌ�&D]����f	���i\����(v�9������m�X	�[�T�V�?=�A�fZ�/�/F=�^\��(�~ņD�T8���ϣ���4�~���ż∔ܤ7:�U����<!ʘ���1�oe�.�N(P"NC���"�����>�L(Y0�k�Lm���LTiQ��*$R�2��ٝ�z���᠉�#|+ ��]�7���Ƹ{w�u��U"�Y��?S 2&1�7�³�a8d�� +�$��y'�ZV�{S�g��%\A���c�M"�Ti&�FUD\*@	ݦ"�ئ#���@��#!^=��\��W=\�ٴg$����6-S-�x�
��W��s�لl޳�L?�nvz�C�T�T�g�1��&e�&/���$!_X�E'(��kdEm�3������k���zS�c���\x�Q*P� ���+v�M`�Lpo{�uV<���;�&B�+Q�o����ʜ�jgH�*�"{v���2�AJ��h@T��Xܡ��֟"䞟�~7��|WR?�+�� ����ޖ����/�~���`�s�+�¡�;{��t��y���P
�<���ߞ�obuFջ5��pt��O�L,���hu����lCJ��|2��ٮ��3ښe���`������V0���/�.^���tx���up�O_��@m6Z�c�ɓ��]L$A�/�AH�.�#j�gl9J��Qʀ�A��s��l��_T�]�h	�`��'�'F����!�H��|�Q�~�Ç�Ъ'X/�<�;+�Ӊ|`��9�~~ΌE4��o�>1`��L�`3���錩����|�$^A�d\��V��:�ȗ��Z���� ?>Q�v27��a��egf��w��M��͍� �����^y�ؤ�}~��n�39&E-��=�
BU���j���AO	h�c�,��1�$����g�7���ۖ�,�U�4��.�oT���Ŷc)��s=F��	!��=�k�L��Ǹ���!�9���9�r�F�qy�͟����z���Z_S�b7
�����~Xf*�3��W�9/])X��t�Mf3�KnR��6�&�'��q=-L`5���3�p�Ք��J�ή>�˖���_;��XN�:�wm�J��}
2��S�OXf1�� �q�A�-j�Br�_�> ��'�%��
 �͝B�#i� �Z����q�v�I��i~��~^&�����@;�z��oԼ~���������}5���nёf�� ��,	��Z� `���U��H3�e�ղD��n5�X�j&v��E�=�H<!����v�~-D(=���z�|F���ߦ�~�� 'D��nS���uKDL��j���9�
N�k{+/"7%X�XsM(*�W�\��lW3&( at�8����s�FL0�_۹��AV}W�^��^)rR�,D�Mo�6=ﶯn���\�B^�R�$a E8��-Ԩrڭ�A�vU����}��l;��mo�5�G�I�̄&czm�%�gY<�g�q���|㞄O2�_�Z�6�q!���Bt3r�7� `��5�g��L��6����	�Z���2خi�� �AL� �ڽ��Sєzq��)��ސG{�Gl$6����l�a���YD
��T�t<x"�����\��B���S ~�x�i2�D s��oq
������(�������a��O:�����m��˸�R\������u���J�5�xZ<ùS�U̾�|{R�ZŷT#����΁_��{{��ﻐ��w���}�U��Mf^�q`���0�3-�?1��e

�
�%4O���(f�b�-���L����r�9�-��>�I,��3�)Hsp��#�sP��2ҹ���ţP������QG�?D��0B<��Ӈ�<ck��t���`���\>���D�C-v��^��'t	9��ե�1<��ח���Y�ȯ�� HvtZ�R�G^FY"ԤM�tf �n�ӯ����PX���9�ॢݚ/�~����]/��= �2�%�e �qm�l ��:1|��]A�!�JacM��Đ�(�$N+��}��
&��⁸V÷kC1����?'#�*6,���1�u��/���G/��p�+mM��C�3f��3������Q���ڋ_��x<�ӕ�cOG�0ý  ���N�R�c@-gr��h�JΥ�)ǁ#Z;�).k�}�%C�=z�l�;؃J����&i�+�JjFHx)���՞g��YV�G�Y�yUVj3la�t�%�1��.�f5�x�xΨI�A�#~7q��1� �U}�n��2&����ٍڼ9�~�)�ޭ=H�:R	ٮLR�0���F������FN^�M�z�n3 7o�����C�y+&�ru���s<�_2�B&��v�VVbn%��e�l�ƴ�~O?)m��&��`���1%�qLܸ�,1���ouu\�7F9YYsYb_w��&)4�7A��;Z.I} Q�T�O/�O@�n~B;����v��C���	����F�����̠��p.{A���<��t�뻓Q�e���1R�	�d=6�e��7��  W����I���p5篼`l�Q3��$9���/��lG���<�t4�S8�c4��?.�\ei wk\���1=�xIag�����b�.�?�˥��D��G����5�-n`EjAFw,�;���Ȥ�?xn4�[�/{��}Y���}U4���Mkx`����j�\a�:�昕�<:�+�00�*���K�/(I̥���Ǣ�A�c+${%���D����~D���p�B����>R�b��}��3����E@��_�43_�D9�;mxit��j����H5>)�8�����~0����ZQ�_���K%A<0
�Gۼ!='>'Wj��6~�|�r�
��Rl�v��.X��h���[sa9�t,jis�}TF��8�%nߢRuSNYi�m�z�h����{BByB���b��B䪡2��@��u�i�)n���������I��Sq�	�mϝ-��s[[��p�>	�4��g��#��1�$e��@�`�	-Ħ&����7�hF0FcФ#�"����d�:���*���A�?�%t���/M{6��F��7�,�bnUc�1�"��~���L$��t
�hɰq��D��qo8f��>f�-�l?2|��`��[�q�oUK����GL�e�\��\3�`���(FIfo�p��k	�5'a[�hn��g�#��;��@O����[�	�n΁�S�0S���SG�v޻G�p��9�U'�ׂù��Vq��:Y���2~�G�q�s��$�Q+Y�?�h��=��8٘Ͽ��]2XN]�a�7pg�p�M��l���}bI���2�1�=��_��y�t=�m��8�"� �%l��#I���w	 ?#�`�)��1C�uh�ʇ$�����bx��29B)���)~��u}�)�$S�]��+,w�Tkjlm�sao�nf\�� F\έҞ�oؚ�v�3�K�u���~	��\C�(��R�DP����ǋWsD�'hK�.KS[��ݲ-6�n"
嶺�Omqv���yq�&_�᫋l����iÜT�=���J���D�/T�$Q�ThJn�&Є�!ڣ_�Ija��;���Mo���39[�W�a����r�ě��88�h����)�5��(-��SS���O�R����nTF�&�R��ŵ�۷w�@���<�V�j�HW���}lf�����2�h�dQ��z4p!;g��%l�?���ȉ�R�|jC�Mf�������c���Y���
���v}`���jw�Z����<���+��!iX��0��ӟ����5� ���1�x�q�
�ɞ��ٷq��\���-�u����un�l�ږ���>l:"̤�H�S���.��72�!�e8g��&�{�5�2{u"&a��ϩ��Ov�[�&�����]�ҀP5�6�Ju�q<;`!m�x�q��	_]���B���|, .kMv��-��>YO�e�n#�#�Z��q��p&)�^�����A��I�6�k3m�>_�O�$�dS?�h}����M�釔	&y���:|\�οw�GĬ3��f:]��ȇ��C�U����?��M0�A�[�ɦ�B(%�3z��ȓ�c�:�v�V����s5ȩ�j٩���S�"��>��YJD)ո]\ڳ	��5�f\�||q���/��@��jM�p�)	���(����μֶb�w�<�W�i��2L�]]��|]��DH&nM-}A��k�����\�n��-��j*�؝�NmTH�fap��`�v�>VJՖ~��� ���i.�Y����^��$�?(.��M�C��Ir��-�W�-d�Kd����@��~�/l��y^߿>��f��2�1 +E��|'O��-ț��ط#�h��_ղ_������p�{ۺ/-'Mmk<��E�>�?��Ʌu�����e"{B�&~�=���5�&��a�%1�_�����B��:|�k�T�|�����ֱ@�w�s�a�V�>�"��ǲJ(��ա�1�/�D}f_g'�b^�|2w�tL�K���L6Ҧ�w$P��&�u�F�WH�ەK�$�����������]R��@��6������ܦ�>9&{2�k�v�7�"'L6^�&�C����W3��H�W�G%�g�!%�����'�/>e3w�i�kA$j�QT�!d8��t�y}�����6�����+يcb����d��vaN��o�>�q�����,����})�[�v/r����#�FYF0��2����i�!�"��u�֪3+����L�z\]HyʑS�f��؟�_U�\�	��!���.���5�F<��.���:X%����Y"S�חl�C�]�lϞ����v�k,�������ͻ_�����a�pj�Aa��xN�6L��m�t /#H><�7�C���5p��J[�I,��H���$��Oo�"7d����\�v��ѱh�]�������2�M�~�^�PR�܊L5�����N��*�BMs���F�����Ֆ��-f�'��|6�wO>��5!oE7�|�}�&�o\�ѥ8r�gY�f���,�
�˛R)�y��g��m��ǳ�3�UΌ�5�m('g(��{.�Yj^e@�R8��x�_b}��%������$�Ğ!MżF���)���o�
�� �;�!�#�+֓tAo �<���^�
������Ɓ\���z+��H*q�m�>�u�\6��>D��M1�U�mSq�Lk�C��I(v�mီ�Ap����2�z8̰1�Y����%�pk�L�ly���ᤐSȲH���[���G{�AE���k�Ƶe^˾/]��ǥor�f+�>�"Ȣ��%�]o�H�!B�Z&�v*���������U�8U��O��z�Y�1�ֳ_��r��Q#XF���?�V�	�xٷ=7]�=D������Uq�G�q� l�����?4Pk�p~uyYRl�����ʶF�<��D/kr��CO�ɣ���ڸ��ޙd-�KZ^7��f0���,�e���ÎV�� ���9��>$�X�ɳ1�����p���#�R���qL<i��m��/��wiɲ0�6�jt�n�j����]I��2����:j��m��G�&Q�E*�Z���""��f�c5C7��q���7.�=��Fl�x��"��҅$k�|Ǫ�g�&�%�������}����
k~T�$WT�B�.O�3E�5�����R8th��.a[
2�럇!y�e�)_��a<Z�01$�����	��6��4`&u�!ʀ�1X򽙅�
��G8��jFH�K׏�w(�����ѺH��T����gw��fuhrx���Ӕ�%���}?\ f���פ%������Rƾ���lAja��L`_a	�Y�Ѯ͢}b�:�;���[�ul�<P���K��3��[;�iN�^A?�E�M:���bB+, `?l�yYbO'm�~��(y߄�ط�'Ug� �}J��|���tCF�cK�M��0�(��i>KQI����X�7R�≝7���H3�$��M<���q�-P��Ѷ��HR�Q0��!�F���+�V]��]�vԈk]�����w��3�H�u8EX����I�Up���Y���]y�ߛ���eJd��_U�n"C�MrjP �V����B��d����<�!C�"6Ò�,Fai0�0?�T�;AB��؅��9Wo�K����'����)Sv�kb���L��qt7\^Ȳͷ�����(sۗ��ʗ��_C�kB�W��01�ә�������
�ÃԹ�\}�*-�l��X��`�"��-���P�sԡ
�m�Y1��0������|�Ί�9��z�3_�/�F�>0�4�7�t�[����%���C��c�1�V���]FUk��^TAHaO^S�P�* r$i���h#U!'{���y7���W����q�J������c��C��t��q�_���g��cUAC�)�=�J)3��J�X���3W5�̂4<�� M$H����Ԏ�M�ֹ�����[�k����+���]��R�5u�L*��f"�q�󲰽��`Ɋ�a��zSX��É���� eT{=�b�&�[6��B.��qm�O�.�[֣fJ�kDȸG�ݝ��	N7�K��wJ2�;�P�!�"V���|�>re4�8�P�F�� �����\,��YZ7*�!PU�#`�{�xb�<	K�xs��h��5$�Ǿ�J��|^:��I�,�|��!�@�m������=�A+��K��'}��
AI�t��$táQ_�b��q�F�`�B_�] ��!�������Y;��uzItG��(������jK.�����X�7����99:�yBY�Y�Q���%�+�Z���ރ�բ�J��.�-��{~f.Q�j���P_E5��V2�Q|{5�/�����1����a�VbRAh*��l㪳�J��i�,G
�h�$\�n'���?*�cOZwi�<�ɮ���_b������ �4���y�A6�sX�����ŭ����0��_-�&y����=b����K�L��nۺ����l@$�qm���d&p٣ww^��6�� ��}�zz*�w�.��QR�h�z��I��h1�}��1F1�Х����o	��-�i_�.E�apҊ��8%�wS�?�0 �̨>����v� +�	o_�mL6�I�Đ�����r�&�j�Dr
��_E���%ve�ܺ�����[� [{��i�.�ڣ�p8OLU+lc��N�q�o)We��/w��|�/Ѡ��Pͷ"G��.��Ĩ�ߐڇEg?5�~Ŝ!�I��S*��g�)��4HN/z[�2A\���V�PR�b�/����w���nr�\X��4����RW��&�����^|���C%�G��>��W�Ua�{����j2:������63h�/�R!�5�!�/��Q�s~�}��d�w�2<=s��(6i����I�5mJJ���E��4���	I���Gӝ+n�\ī���􍝋�o4��]����Z��r&�����T
��6�'�'�=O%u$t�������@q�r���k-99���o�7�m��G6���7^�T������:�<o�M�]��Ry��$f�%3愵K�7�A!��)�A�	zg�f��z�ᶨ���.�C�x����9��)ص$��x�����EB��P��uTJQ�~��El=��Ҫ!r1�ǪH(�B�y�Yi�g�0~�J:u6����.�Ɇ��vh��}n��>�L�Q����ƪ/��-,2��}�C4=�U
 �೿���F/�Cd�Oj�&��T\��n�&�Gr���6�H�.�}�Ô�Kϯ��f_>���������bI=1��lo��*��>f��_�Y`�]"��0�{���,��39�5�i�M�f�u5S]���S�Ԃz�r���@�&��0|�vwl] R��TW�h��������2;��%xNbe\�n�B�����+�ѿΞ����Susk_�9z#D�L���1��� �+��m�iu��%���4� �'���)a�q�~ה�S�	]z_��ܨ�[_�T����`�"`��b_���v���V�>,���#CĔ� ����\pO ��X����p,�	V���գ��v�Uj�����a�7��������ag��� l2�M
h����
[��K��1ŷ���r���]��[�@�4mB�}Pފ�=U�W�,�U�w�ۤN-T��?+4吽0?Q���Zv#��Ӳ� �Ķ��]vOT{�,'M�ۇ]�`\��ŤF�'�-z���Ȥz�(b0B��HZ���E�u��6y~8r)��_i�Y�9�)2�R[j�5��#"�૴Z�U��4&����r�G��`����\/EG_��|N2�*���.����$hL�̰��a�1��T]�Kc��Ɖz��'谺j
�Y �B�w8�Hi_?���
W�^_2/���.�V|���Za�y���Ee=at͙�Wo�V�$���o�Aϗ,�E,��0���0n&N"��V�ftѪv�?sZ�PS���	�i��yj���Գ&�������T����O�\
�2��'��y�@�^[K���:�O��-�Z-Mߙ؉:՟A9Nz�7�sE> �¦��� )�<�ʮF�faP ��
#-�R�����H�8Q�� .���z�Q��ή;XHl�=|y0���hr�]�RmJ��Z$6A7~�ߠ��X�-�)��p��W���C5C�O�` F�B~��֗±~�Ϫ�|v�%?��p���D��ESF�{e_����|�c�����&@�W:�"�$3E�L���=C�G��d��H���%ύ�[_7=��g�	�mhu�K�����/��% �3Th���d���uԶ�O����U��D%w�K������R�us�����=�����S������p��~���$=e����C�+S�\ >_�r1Y$�5�&�����y�\�����`�:A�ת�H�&7�r��A0��'r��־ؿ���cD�f�F]C�b����r��ި��S(�|���t���7B�=U� s��g���:GC�(G�/N���@"P�	�@���r�bBUy�ݰ����ƣ�m�m�/72%�&Q�������u:jG=����Ġ�KՇ�u!lc�I:bf�[���)r��0�0�8~9���la���۝P�1�����X�/�ȼ���3�F�;��~�9�V�����6��#�����+���2�.Z߰�3+��
��{c�
��xW��%�FKW	Ta�s���B��VI���m�9C����̫�����v�D�ڕ�{d=��g}�k��P�������P(�}0��iU9c�Β	���# ~f�����@ w��E�r ~�P�:ybJ�iB����\��Bdע��5��l�
=� v���t;�{���U�;����X��s�\��r���PןK���x����e��8����
���L i/��Ip�;Z�_D@o