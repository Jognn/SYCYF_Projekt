��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&��n?��1ů��> K�-� �&�T�Ek/ֆ�\�놭5�DꢘP���+L+X�4��J��#�0�8���������l��jT��+�(���������6�MC!D�;�m�퓊D@v_p��䙋ⲝ��C_�6�Ռ��#�� ���	RD�4D��畓7���vn�H���0���fX����4 �CS�C`{��;�L����li��� y+����FD�p"��]���y��R��K�({� .؜M�������	^5���ɋ��&���&�@*���
e�� �t+���
_6��O<��7f�M��u���m(MrN����z�jL���@T`��M3��c�uQ�Y���%�dD���,�~^���y@Ga��(����C����	��G�86�S$��ɳT�ز8���:r��/y�[ݦڍ#A�����i�&<nU��<[5)�Z�-Ĭv���0t���d���"_���:�'-��d��*��q����_d�y�N-��~";#��������Y��؆���	6ZJnԷW��έ$Y�K�?�4���L�w�Wmiɶ��Y�?jx#*�i���F�m�E����O6T>]i�_�9;�!(��kH7�OS��_��[-M�((��lO�s�$�g�x7`��ZV�E���F��,9�j	@���]}<�ahb5~ãdl&I^�	v����-�@�@���	��!��d��`j[Q��� r��;f�i�.�m+UH7��/OV��c��������l��i��M��*'��?���G� SK�M��H?�מqT'J,!A�h���'� D��G�T�>��tw�ܻ��l.pRu\7�V-�T�V���CS@�ewf���H�*�cwl�H��ϋ��#�`IY�k����_��U�A#���z\�yz�~�cٽ�bl����S�&+s#�V��%��ӧ'A�N��qT�7a�t��$d��]sH8�G�?����i��i6�ˋKl<�O/���	w�C��:�D��]�l9�ތ�G6���Ccyg9m��<%���o�m:|0�\)!�)�2�*�y�e�M��%����� w�Y�.���,���E�ٗ��N�*��O�zP�i8:³��v�\ݏ*�P�?���`�l��F-U=7�g���w��ȩ��$���"5��!������{Kh��������k�$V,[No�"a�K��H��c&W���Xu3ѳ����i�uI(of���p4<t�Xzf��4p-h��,����<��W%P�)�������c�%w]������"� �ۭ��9�[�Z_���K���N��� �{����Z�@���k}]�s�yR��݋}�k���/���7�&�<�V�0��dG�z}af��5#8��N1�M ��Tl}JĖ�B�	�}E�}�A�	K����D'�R�g��=	������+a������%s,^m�����Ԝ>�m�����?��/ ��#]>؊uN�\���0}�ڇ�T���cj~9�I/g�~0��1���'`p�4��w�:�)�W�M�^�p�r8�^�XO�>j�̫h��BZ�T:�x��z����p<xͿ`����u%�����HM��@\�(��'��b�#d�O��b�i� �SY�L�Z
�=,��H�G�tu�>��^<�Hv��o�z�@�(&\����F��Fq� s�SW�Gv��/������bE���9b�g3D
�'��}d��s�3�KZ�+J��#ӎ���<0}����@A�k%߽����ș39���G�Zx�D�\i�i��6g�i	���hpw:Pl����kϞdKl���<�aK�'�r��̯'��!1�K�cZ��`78��"2�P;
_��i�~��t���p�.A����#�,������V�Vj�+:(���,(�ajƯQ�P�L �w�9m�l�M�+L������Vh@:*�ث0�8ھ�,7�4G�7>GJ
�ǃ&u[��o��]u��(P�Ҫf@[�ܠ�Hq�v-�� ��?���@\�0^Do�s�><�]�{oZ|���}�
�{�Op���ɖy*�Ҧ1jk�xJj�����j?��6pG���u3���w�>2���B]L0�vBP��h�J�OrԒB���%�c�^�JCw++<YTBs<�	kY͖��&x�o�2B�U,y��]p�:k�1����](7X*Oeᆇb�T�AH\��N���\�K��R2`u������st�'�//�8r��+�@�×�?^�/D���6Oxh"���üQy��?`/��"�����"#� �Ū���������  )����8��pD�N�&%*�R>��e��N�J���|e1v����JR��)�*��� �30�Q�4V���/W���G8�Yўt����H�����d@��ͮeIe��U�"�,��L�'��ꓰڇɢ�N��s��b�~P#ʋS��y"��2�M�W���}z.k�i�y�q��M�Nϥr]�(�A�}��`����? �|����(���J������<� n����(��<�na`�sO�F+���q�nL�t+9@u�� ��'��T^F�O�c�N�F%E6`zb�gnA�_�"
���4tq�����ܹV�B՜,,Gi��ӑ#��wZv�]� O�]Y>��W���8��Aw ~�܂���TWv�a�:K�7<x����=@�ֳ����s�W�9@-iU`_Q�D͏.	�I��-Fh���h^���X�Uva�M�=�l�jY�|�d8֖��t>�?O0)�."���j9��$cH� ����v��? ��LO�i��t��X!]QX{t2��K��p��W�&���VL����(��񝪟����PTB��PD�$u�*���+h�P�;�B֎8ԩ�}������l�0ˡ��������v��+�\�3ѽ9*�N	�+i���2�a���2*��$)�X��F����!T�g�Y>���"$�hc��%�{,�i~��d�}�4�T&����|����o��6ȏ���gl᪑�ضPW	h͗�J�
M�vx�*N�CN�	z�� �1��а�W��{V�a������(κ�٩g�p��s�>�*a��o���}½)�!a��[���)k��[Ͱ?Llo��C�d����iU�u����`�0���X7<�Zu�S�mA�C ��� ��܂���.:ak�i�lV��7�U��x_=��f�����{?�l)�kʄߢ�����}޺i�S
G �jO��7}�W7@�^L�1���k�fV��.�S��ٔ�2CWNE�-[��w����7���yO�<��q�A#֟}�#2�<^6ɓ�~�~צ����.�l��
	�fb�5��L�<tq�-f�k렄� X���<���R�ii2lhr�9RyV0��Ǵ%�8ه���� ��2���n��m����AC�$K���VL� #��l�q��&����K$ڇ�dz�1�.bo���`�H�t�n��Nc �Ȕ�)�w(nqK�sI
aܣv��J�CR��B����>	6g%���.�;�5m�~"��Pj0����nDI	�me�~��]���@֎���n&�߁����q�Ь[}��o�<,�e�zg����*�TU���w�^���z}u'=e�,H�ߜ�5se�gS�Х! G ��Şhy��=4�ϼj�?�&}ef�����a�#s�H�I�D���%ZAx	�L�8XDT�$ ��Kof���H:|�,�D'�+ �I��oq)��^+>��1O���spX����G�(���G|��;��POMI	�w�V�T�QU9~18�����vE�t��g���R�h6�Z:�� �qo֬B=we�5����t���`;��3����'B�u�@ߛ � ����od^x���g[ck
�jc�I�t��>�(ٻ�i�/�_)JT��6�a���n�g�^rEX�i7��<�c�ִf� �����W�y�vE�e�����߽��kT6�i��9ŏ�#�>�i�r8�$|ܸU�T8���{_����l+�xg�����^߂�*10�K�1k��
���Ԛ|@k"��)�݆J]n�U#����0D5m�����NǊ����՞��]�� �U�7��/$U�-#�7����̖"[�Us%4�t��Plźqh�x�fΥP�˃>���X
�`l~���f�3�d���6���e�3`L�#+���Zov$J�צ��B�\���x��^�3�L�h�L�e�y�
�Q�}!;^� Ũ����,H2*�"=����s��Y��<qI��]����&��%4����ڌ��|�]zB
�P�,T('����".�׋�y���b����m-mԀ�|<���9C���6�chڱ��n�{ޫ!��I�<[�8+��w�B�j2�s����4}���r�t�Y
���qY(E&.�,r���И�!1f�2B�ծr�ûź���]�]eVt�~����_g`�`d�Z�<<��XԤ<�mf�J�g��2������O6�v@<�Q��P܍.��s�|8��$Ύ�Js�^�tZ�P����+5�\H��
�z5���eK�Q��I�ᐺO����)�<r���|���5�䎛�[�߾�lv�gkm�YC~�R+-ײ��Ч	���[b<7�z-9L:�c9�(����K�t��/����B]Y� '�Tl�눪Y�;[J�!Y�i0/�
����G��zh��J�k\7��z�K8ۂ�B��a����������	�m�0��̤;��2N��G/?��]p:���Qx��y;���N��@g�LI(��H�ߊh�F��N:(L�oȯ��[�<{�-J���3v��Tw�7U�Vp������, hD@�N�?�?q�6��QM����yܐ�3r}�L�pi���	��0 ��� ?���$^�#�O�a�����>�=֧�J����S��GPL���|��ʎ��!�:^	��/^��u0���9p�&�A��4��0�����(��7}��s[���(J�9�����K�@X�.�p�st��td}�U�+�<|��Z�o���������������g���ioQ���9��SM��c\��
6��#��!l�G-��i����eʎVL6)b����Zz� #��J��x{�Z��̦�7HG���~��؏@�9��J����`B�������X��vk7��8�e��K���F���h�����ju`!0-Bj��s��[�wRiZ�Qqɒ�p�2E����@��L�����S���{�T\<'�Gc��e�AlWv�'W�t�8�\ݗ��\b�����mp㔵9�k,1f�yE��l+=���6�Zz���� Ѡ��l]��%'J�$��+@�^2��������>��/��Ų�]�Z��e���P.����Cx����Ӵ��{ɂ�J� b;��J��Hd ��vC!a�_� }��xV�VW>h�Ի���#u�LQ\<�Ϩ-дÇ�n���l��Y?d�-4+l�rF���դhl#���L���Ɓ�8 ϖ+�K���*0�մ