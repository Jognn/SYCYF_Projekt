��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&��n?��1ů��> K�-� �&�T�Ek/ֆ�\�놭5�DꢘP���+L+X�4��J��#�0�8���������l��jT��+�(���������6�MC!D�;�m�퓊D@v_p��䙋ⲝ��C_�6�Ռ��#�� ���	RD�4D��畓7���vn�H���0���fX����4 �CS�C`{��;�L����li��� y+����FD�p"��]���y��R��K�({� .؜M�������	^5���ɋ��&���&�@*���
e�� �t+���
_6��O<��7f�M��u���m(MrN����z�jL���@T`��M3��c�uQ�Y���%�dD���,�~^���y@Ga��(����C����	��G�86�S$��ɳT�ز8���:r��/y�[ݦڍ#A�����i�&<nU��<[5)�Z�-Ĭv���0t���d���"_���:�'-��d��*��q����_d�y�N-��~";#��������Y��؆���	6ZJnԷW��έ$Y�K�?�4���L�w�Wmiɶ��Y�?jx#*�i���F�m�E����O6T>]i�_�9;�!(��kH7�OS��_��[-M�((��lO�s�$�g�x7`��ZV�E���F��,9�j	@���]}<�ahb5~ãdl&I^�	v����-�@�@���	��!��d��`j[Q��� r��;f�i�.�m+UH7��/OV��c��������l��i��M��*'��?���G� SK�M��H?�מqT'J,!A�h���'� D��G�T�>��tw�ܻ��l.pRu\7�V-�T�V���CS@�ewf���H�*�cwl�H��ϋ��#�`IY�k����_��U�A#���z\�yz�~�cٽ�bl����S�&+s#�V��%��ӧ'A�N��qT�7a�t��$d��]sH8�G�?����i��i6�ˋKl<�O/���	w�C��:�D��]�l9�ތ�G6���Ccyg9m��<%���o�m:|0�\)!�)�2�*�y�e�M��%����� w�Y�.���,���E�ٗ��N�*��O�zP�i8:³��v�\ݏ*�P�?���`�l��F-U=7�g���w��ȩ��$���"5��!������{Kh��������k�$V,[No�"a�K��H��c&W���Xu3ѳ����i�uI(of���p4<t�Xzf��4p-h��,����<��W%P�)�������c�%w]������"� �ۭ��9�[�Z_���K���N��� �{����Z�@���k}]�s�yR��݋}�k���/���7�&�<�V�0��dG�z}af��5#8��N1�M ��Tl}JĖ�B�	�}E�}�A�	K����D'�R�g��=	������+a������%s,^m�����Ԝ>�m�����?��/ ��#]>؊uN�\���0}�ڇ�T���cj~9�I/g�~0��1���'`p�4��w�:�)�W�M�^�p�r8�^�XO�>j�̫h��BZ�T:�x��z����q���r�q��_:h�q����Y�}��]P������E�
����
	qZR��+������XR9߲熌�������o�g�{�¡����7*3�{�ԉ󯠎�ӼW�������\�	G�-Kٚy�����V��x
�̒�}������h�Yڵh.�W�Hy�)�6A��6
�J¸�������MPU�l��Y�9�LE�­�`����+���eo's��O�KZ��\��:^�u�e�FKE��m�y�����m8�^�^M��zfJ�QP��'��d�d-�]��U�e���4�B{���y&�Y��Eu0��y��r}�!H�2�-v�����<y;\�q��j��O��Q���P�퇑:�Yge/��%�ׄ՚���kS.,~��c ��.�d� ��9�y��y�Z~�o\�!�(.���=�Ă��J	�h��ؔu�ɣO��o����XɺA �Y�j���!�lZ?�bƃ�8��N��r;n��z"�
y�bI�1��q�(\�\����$���_u;}|x�8�eo��Z}�븎�f��P�]��9Dw�n7���i61�~'g�՜���[�6MPN�t��yb�J �X�t��f���:�;�&$�|.�X����F;J�Y�sZ�e�#]o0���L�$�4{mqپ]�K	�×b�(�l[�����o�
˦��e��������%4����9:�UCHZ�/�����=x�'WƂ��;s��#����p���s��{K33��\�l���3�߮?ke�c�k8SC�4N��$��V����4XտTsc�c����s�?�����cb�a�"(��u&����<�E���r�q�D�Fv"��g1xl� �j1�J�.�{�9�I�����R��b�(��pN�G���������s��a�W�&8ht�� ���H�����OF��Q�EJ���f `�9z�mOG�(A�5~�:R��h�,��!�}��p\p���Y4r*��P�yOB{Z��������J����R�2{��Upz'����r�!�ȝGK�4g�� $J}�J��ڜlW`EԤ���Z��y�`$��Q�W�c?o�$.�հ��]�n���E��A�3����$�th�
<��L�-��tKz�hHP�ltD��?I:�/��p�qZㄅ�S�-��^j���{}is�����:	����nJ�{�E���|@�&��]<��	2�`�g�Ӥ�N�&���Sᇢw�cl�m
��"�1%.\����åN�\��Y]1২���U���\N�/�vB��d���J�M�fR�o���.�}x�a�I�6�L�-
��]`}�KQ �+lS#��c�Y0�?W�"r��/�
p-'�Mٙ�E��/��ōW�
o�Y�1+
�Ϩ�&�-+/;e��>�o���b�p�M��f�9d�](a��e����\'���R�]�tBa�w�dE^L�����s��<�*�C�s1����aj�x=�Vԏf�_��|TKV��A"�9�o�W��� ���3B��G��RK%y���:�ѝ�Y,�0�[���@']d�0�]�Ֆ�7��TD:�׮[���7��=��0D)�l�h��葎6��#��_��Jg�9| ŕ7/2i'�<(����� D!F������&����JT2�<�������ͫx�������x���Z5�GBRћ��	�\�')a����3l���[�n<E�x��~�5�����=��JD�+SO��[>�P<v� �-�q uC�����Y�b�/)�-�0!(� n]4�/hg��2f>����7�b۰�X-<��*��6e�:g&㣪&j����eM��
���ke�D�u�e��M!/�X��_P���T�W�~Dﶫ�U��t+���� t�t��Q�6��('�a �	/��r"�㩗WF�.��?����B~jX�;�-\M��������i�Fv��M�R`^�i��^���'�Pƈ����e����E�doo-E?��S�e��tP&*�V��Vܳ�x�\i�f�!<.���4����%|1!�r6Ȯ.�ͧIg/���n�ڑ�e K��a)H D�ڗ[�5&�m�M  r?�?`�A>{�H߶�p�hގ3��J �����e=	�aцG�f,Ͱ�\���F��N�{��,�[Oǚ�PZ�XR�p1#�lE�/QK8�;�@쐛:��b9>ڠraL�c�$_�2$<�=���z&�!�0
W�!(��W�t�((Q�no(!�(F��o�Ϛ�]�R�9t��zi���?�尳L�!$b�Qڥ��1���I2��Ki;�5|�����:�>:�s�m�0(aF��G�0���׌6lܞ�U��&T\ 6�G���<�6<��omH2��#Y���@]mL�~J$����AA��0ы!�Ù�0�k!�� /�^*3�T:戫E�?I�Z��ʀK��Iz	�N/��*���&Y���b��]�욈���gc%��>l�Y��!|���S���z+���[�ٵ.R�"�s�q�z�<�r;&�� ɃD��c�e9�+�v�:�O���s��9�ˋ��'��ю_�r�OE,Е��K�����;A+u(f��ݯ����ao�7#C���q�+��{�*G}?|R��uu �d�Y-�q�^�K&�v�?Ɨ[
�e��Ud�.qk��rCr:?ث٩�*N��U����w),�2$����ʤ�6�s�����0t����^P��,�����"�]�l�5C}2y2=�J��S���DX��s��`��AF��,g��(D��gXU#�����m��^�ϯ�BEG{�4oY���u�$�-b�0	��]����9=Х-
d< ���幆K㙗�eY�E�~��V7���,7�S�Ci��T�غw��X��cv~ys�i�
��`^L�.�3���}���~��p�p_�F1T/*�V�╠����	��fK۵@�W��6�e^wޗe�o�epZ���;�P�us�^Jz9C��C��~��K�s���}Z�y��:�.b�-|���Y�:1q�����O����g���&�Q��UFz�o��l�@��@�{,�M�|`+{���^1��N���S�Hޑ��� 3�}(��9�=�[0d�-z3dD*s��}���6B��h~�Y����rn��'Bl�q`g��Z5����o;���N2�R��V���B��1��&��A�̀��5:�֤����&r��O֎[q8݃R�������J���HSjQVK�q�d����5�+��$JƸ��Lsٞ�C����m���g�v�±\�.S�s�Z	4Q����n:��M��u@:�{�>��{o��������>?0��a�^<�{PrM)�Vi ��|j���6�r,���=�7)���UQ^��)ئte��?Dڼ�_M�N�������.����;�G���YguʸI�_���S|j�|$�TCoS�8���.��C��lϬK���[V/:Q;kU�k�w�������s��qa�D���To/���6�._���~�3!��b��c�O�a�����FR�������-K;�y3��w��q1k�%��'�X�:A��}�v9B�`1.q.Z^'pf�f����N����MXJEK�e���e�8�PV���Ի�c~p,�)�	��
G��i���w��H�ᚫS����8�=s\��:�^Haa��_��#Ӂ�HO�	��`yCgX)��犫��ÿ�w�0�M�3�'��j?P��ד�*�)v�r2r뚞������9-k�D�<H��O��@�X�U��Q}��8���T0t`Ty(�L��:Z���Q[D���>�Il�[���Z8"{������Ѩߪ/XL6���Y=m+F/���M�90w5z�l(cTwy��N��K��b�U%z�1e�뗛w=�fsН��b�/q���o"(ѝ�. ���> ��_PtoR0��Ďv%%� [,f49�e��1�O��7t=ER�{f��F�� c����a���<������\�^!�׽��M�p��;���E�-B#�LK��)KE���fH���~U���bpӨ�ޒsu2Cȋ��_$.p�m�%�A���̫����w ��d(ё�,������"B,�Y�K��t�%�k�R�<Q����2P${>2O�_���%9JG=*����1m�	�c�V�����V*��/�m!T!�J#��#Rg焮���� c�l�<�Ȉ�#�0Ę/#if:���R���R������9"�^�D�V`~��*�8O�A��PR&H�9C+P�+G*���5 �v��M��U��ſ�'���R�W3��UY,D�r7��5���g��Ox|p��Hzf�Y{�IC���<wf��&yb����U��c��@U5��l�()�1tu�"���(}ԑ�a��@�������}O�gR���p�Oxd��¯��g)[ޏ�p��~G|�%��Kh,�I�8x��	a�Ł�~-�7��[jxq5aӏǫs)�|\���|��zI�
$ɜj\�|��67��)3�q��8������=&��Ŀt)�{!p1�m�q�i_Xp�vFD��g�D�F:�B*qjhb��*^h�_E��-�/|���	���#L�sz�E���ky��񚭆>>����j���9շ����sk�5�=���#߇R����X�t���X"�o�dm�]̿AxYf�b���6�"aҶ�i��4�_�_ʜ�}xƉ7}�����*�U~�������d�(��#�QId(����+eQe�5����ek�P���?�kN~�I�L��]���0��-��܆h���߄��a"g��Nm��SLڤ������26��#�_�|��C*�ܷ�wE�I��*� d�I�ܐ,��n��t�#�m�1`n�al�z/QJ9 넽�^ck�س?����'A�R�X'C�j��/:�iJ*��Ϳ:R�6/�V7�T�G#���x~���!�o��WȒ|�(�j��[��d7;K���bk]=9Ȝ��N��� �rԴg��H�P�@��&j
8�ů4����8�/�4�
~'.�2)��E�'_#ܬ;>HW�B/��[���m�����9�L���h!9��\y���RBMbb4m}	��x�5"��2R�C���ѷS.|#}*_-G�J��H��Ú��,vh'�kܙ�c�wP���@l�-��&ޒAk��3fq;���P��D�ՋH!M�h���N�#�=���M�M�+b���(�*m�7�i�~w_�K��[H鳭���O�4gO�g_%�?9 آ↨xZ�u�j~d�<���}�;Ϲ�H�<�8�*iPi9zl�Ò@����ׇ}b*��-:pKu����{H�Մ� �A>�b�ܓ�s".̏p���_������	�>[)�#e/�J��I��^.b�I�3�]YF1�ۺ�H=e�+��` ~0`jGn�辅_����_���{2�ZƇN�����Ҩ�f���W�Zs(�2�ai�6ĥ9u0[��#�ix"�����P��E$�?��~�N�4�Wr�lՎ3�1��0�Ih���MLGY��XM�ÐN�%26�-E��CϷ� Ľ��o�(7Q\6����>�ھR;�(2���o3
�T!q�THT� #���\�қQ}�iu����ܹ^�80u���iOD��&�l,��iuz��,�+��} 7D��)��b%�+1�� �Sэg��d�Z>�����F��詇��k�lL���a��`q� �WT�vz �_�e�0
���o�|�q�W�������t����P�t~����X�OW�D�Pimr��ӂ�]��%O/d^u�=�@(�k8R3~be��}&�}i�X<j���͂8Y�B����V[�Z>]�)�i#����SH˓�\tv<�T��98GĶۃI�g��Cs�F����Sx�T.}{;L<*���1
��~���0<|JW}�,p^k�&w���Ō�$O�jT���tA6��M;.�B"�&ꂢ$d��/z3ɅC��?�G���s5�4��W�3E\f���8<�C3�M&��:�u(�d�O���R��X���.�c�-�	���>�I�����=c�"ވz���`(j&A�b��׉���U_[�@Z��V�����E���.
F�6��$F'm�6�aߐ~�� �f�%��� �+6���1�o�Z�����Ӷ=�x|�K��x
�k��?b�����]Q�\bT��C�5�Ƽ��.?���c4I1��M=��$�̏��P!�ov/�� �9 ��E�bž��Q�ۦ�aZs�K
�Ei����~~����X0��6�#?�=q�)�k�xu��>�AY�{�J�/�l��DY�ASٜ���h�?-����ww<Y��s��l�J�������������f���4&֋�ť�ڸ�+���hR�鲙^����%�	�o���z�Q����r��'�g�����6/#&\�vdT�a��ծGI�Q��Z�[�M�l7e���f���.��&S���)h���U��YhH+@�<���1��q����t0��T���bx�����!�)�Ea#8SF��j��w�����@룯����J��Ҝ��Ɣ�y8K��֕���[���'7\V"ut[����n,5���y~�����l��f�鳆`�f��Ө@��}���}Y<��{G�S�X�f�u�J����$�Kr)(&�U�1��|��s��J�@KnF $b�ۺV�R$��b�o!t�q�Rkg�z��1 �j�_��ߛD����X��*ʛ�/��B^�ߘt75��T��`��F%H�8�q`^�A�\�"�w���N�H�����G���8���B��b{T9U Ǭ��ٷ��T��-�B$�n�.�%p����Ǆa�db۰%n�r�V����p7�	+��6x5�x&}�����01���Dd�= '��6��u�\m�BÏgJ�0��~�m����-5j�w��0�g��M�;׫��ǯ�ٓx/w��C�2��3���]�k�̅V���%���U�~�۰ �G%1:���U�fn���DK ��{U ^o�U�^E�j�9��<���v���l6�1$RS!������&��bvx��)�S������ R�<��4�UN�"ߜ�{Z�=���Bg�5I�����	�r' R�Y���.����[���ܨ��������jH�0W+%����O���I�����q%J��!��/��0qh���`���0���}���Bx�����z6~���&Nd�� o��5S�6e�+c=lߖc�k��׆�㋎�;�q)⯚W����@҇�AoE�%�B���u(݃�ʨ��i8�P�
�'ʙ3�`�CfP��cg�`]<\�����k��>�u>e~�	���'4��<��jR�q<&�,�jQ��~���J��ƙ�#e������F�4!�;jao��P��xͿM&j����}Y;-C�D-xqmx	V�͕jhĘ�Y��2��P��w���OE�ܔ<���*��Uڟ���{�Rq`��θ�y�����Z;;��l/v�� 2(�Y���ΜI4A!�'0�T��%�~�_Ɉ0��>,2�*��y�=�����^��06r9{�t\��T���ь�p�EK�)t�K3��7ğ`��&[�j�Cg�E[��	����V������	u���LW0ڴy����-y�]ze��R�:S�¨��r.��w�r7&Gn����8��r�v	e�1B�a~�����
����������.y��4�;��N�}�{��J�PH���#��<4N����[�豯>�
u�[�G�o欦,�]�o�wB�� ���at��i�꺞�cj|�����"3�nZ~�h)T92��I��ܘe�U������w�1�Q�h0h �MJ��ߘ3"����|�[��̤���)��ү����A2����&���i�o�_&�TL�;�3��̲�x�� �?�R���;zR�K;l��� L:����9r��d��F��'k�ʃ3�iA:2f��U�s�w�~v�3g!6z\LG��*٬5���R�o#{s���@۔Wo��<|b�N��
��#'sC�dz�&�"dU��%X�w!iݽ����^��1Ć~��)	Ý�� �%��fEv�0�jW�1�WK��i�<�,;��x*�y�>��pƑ��|�3�U��(N<C��]���5vw�������/�d���Ǹ2��T����#��z�3�f$�Q�b���Y�P�m�njܲ���}������`�A�`�wkґ{b�LG�S�Lk��80�U5�ϼ�|��I�t�h�fw_�����˔n����<B�S8���&��b��,׷E�/|�����Af��2۠���Uˎļ� �>jP�C5�v�÷m�2bE'��t��s�S�K�7d�g1��<�!��A���۬r�7w�FK��������=_D͹�̦PK.�K<�I��<jk ������ �kk0=	�W���3�\f��dIs�7�G��P��a	1U(U��Z�"R��˜RM���-f�R�/)�k��>x~& v���s�����;��:H�Lq��u_x]=s�o�'?*��X^v��2Uo��.��G>3MW@,�����Z_͕_shڄ�8F7gX�fcr���+p)0rF��h��Dx����4Z����l n�t�<�O�����׻�2�v�Y|ኩm��EH
U�P�ĉ�@(x�n֍�l�jӵ)u����g�G?��0�:(������w�Y3Rh�9����` T"�W���)�ⵣ������`:��&�gzW'-�`-]�6��'H��~[�x���1ن��~�E�!_��.l��G�<�ޥMO��K��IRJЄV{<�w@�~NC
�������]R'2&1��Hj��3�2 ^rqU�8O@/��)�n+@��?i�/��&��+�ht�4�f�p1r k�1 �i��7�DM*������\��b��2m��,���V4w�{>�N2�3B�֥8��o�j���� ������Ԍ�{;�Y����n���zW|~�Z9/�y�`�Q>��4�)O��4��$vҰ�ؾ{K YeT�p͊fڝI�f����j���bJ�����o����2k��Ę���q� nУ[�QD.��=e5H�z0���r��" ��,7B�R�ZhN,����6���-�)K����Z��l�P��䖮�l���'9]b�6�7&�c�+Q�i�ZƖ����R �����	�u%�Y��<�wo��W���^:�d�(}y�ǝ�e��J^ ���9��}���}�<� ����~ɦ/�g�� � I�� 8�Ӯ�i��ff���uʴ����Q�rO�s �\�R|<̉r��$:��Ȗ%&v���9���ܝ��FJ��n>����w��q����C��(x򽭷y
�"��U����dYF9��HhH��4ҡh�$p�H�Y�S��A1\&�S�q�Y�Z��|�[�[��A�H��K\�o;��?4:-���[kۜ�z~�&�6��띠DU���.T0���B�.�gkp��Q�1�ļ��U�g���t��ΊW��L+�50���+ۋ)�S�Y?�u�I�ϊ{���=<�ӊ�ـӬ����tk��)���TN�Y�n1K��|�T�e�אz�]�i��-�Ш�+b���'&�a�ONΩ��q0n/Դ�m�h[`�̶$i���l|¿S�z!���C�eK��b�]�u���%A|��'i��hl�q��N� �б���e���g�Ev G�H����+����Xh5]�d@m9��}�T�/���!�h��sD��D�1d���M������v=ߌ�Y�N��E���H1QtĄ�#��b	�1W�]"w����woM��M��2ƈB	LE�Q��޾�4��>r�����Q����z$���q�Z���Wqe$BЂB�x�7el��n4 �p�h��R�8�䱯ĥY��U�]�W�)If��G�I
-�u4.0�1�!����4pD_� 8�t�np����p���o�2���J���0>��\繷��!��h�!�rb�����)o��iJ������ĉl�#L��a� Q�����1��d�L��TF
�׭�{���{]�{�--�S��G����0I�E�H;(]B���7`��/�������-m�a4�����7�%�x"��'g��{�8|;���D�R-�WϢ��T�ϝ�`H�.��BrA���?�O�S3F^h����52&�m�T�=�@��a�,���T:�HY��a�٧|޻���D�H����؈��"8��ԋ�����ӕ�L�r�7�����QY,��J�N���X����wͺ�����(���'������	p2���2o�΄� At5-Bt��1Y���A��ꩳQ��/�?Ǒ�x)2���|V��W-~��@�IV�Pf�����h�q�!`��?A9U��(D��ǌo��zc��7`�)k���w�" |)�yO@��iT�ڹY���7�O�糾4����G��4\إ���p�T�_Ja"��Y���5��s�s�Q�}�rX�闟�^�;��*�� �mb���^kt[F�WK%��W�u�2�H�7�Rq��`/��W���;3Ȕ��ĸ�(u�����z@ <OzV�u]��6ґ�r?2����	��.M�*��ټ�Y�䞄���Gy��Zئvce,-�
t�P�t B�Ԥ"{�(A���sq�OM�0���@��S�ߕn.�ef������:K��&:�,�� 	��T'(��ǽb���*��G��!�7@�8�}Y\����u�vygD�}�&iX��s^Q���@����2&����� �m��P��B��O��� �p���h\e����T��l_`PQ�;�����D �H��>��<b"7n��"��s
��mf����`ء�[+��ٿJ<����E�ZS����OϽ����ߡ���P�d��.AC�1�/�r�������}ʧ��E=X��6���1֑�@7�^� ���@Z;�^z�9kk���.j�(��&�F��`�ߔ�)�ö��nL���Á��ڵxW�c��x�0����W�P#XŐr��*
���4߇�p��n���8�����r� w�ӿpIe�sܪ�<�Y�&FAFX����=ﱘ��+v���ByF�j�R�N��f��5�K�����=�NWZ�q�~�/԰z�~Ymh��������J������-��xn�����E^�Q�T8����,U���j��S�"��4H�	�$oa��+6d�e/�H���ޙe���b��G)
X�9'��!5.��{'���4�uC�F2e�!��9��u�=s��q��T��ן�\��}�\MoY q��%�*�sN'�M�@B��ðo0S��Rf%��*�Z=�|�g�	��O5pjO�ݥ���}���+�ۭ��>)9�'�f���i��_���p���_ٖ���T@z|r�_��y�B{D��Ŷ��y�̀�qPOqd(�ǵ�3��4bFD�wO��)6�aa�8�T�u*B�3s����@_�NX�Ŗ��( 1Z��e@˫�'I��	M�Fdg�z�p���{ �,k$����^�����fv����h�'ZB�˹�㮕�
�U8SڪV�L���d�Eϵ�Ͽ��T -�3�,�H}jd�/p~���M�[-��J
UE�A�?����}/E��6<['B�����ϯ�Z��sɬN�#��Y�\��{�4Ed��$�:�de>1L�]��(e�m)��I��/��ؖ�m���b�An�V��~�C�j���姺k�oA{ª���P��I��H��L�`�P:X�*�1|btU\��n1�&�����b>�D�NsD�Y����H���� :n�C�Nƴ��n[��h���t�r��z
C�OL��(�U}���S�]\���o�x�r�TM�#z�.N�J��9�/���!�kJ�>^D,<�&�8譒��(�3"�ͽ���bR�[���#�/SydO�ݞBcZ�jGP]r|����`C��hp̨o�yvc`D6���e�ɶ��_+��PZ�ֻ���[��T�u3�:�<�
Z!s("m�y��w��5F�j�q�����,x��Ln�l�`I�������<�m0����`��"t5�Ii�J���t�hO��,/Y��*�^������W�өF%Uiq�<���n�b���Oj|��z�rpV-�:�u;p�6TڄoT|�g��E`�eѢ�??Vy�Q���l�T��z�$����*㢜k��W�1�M��̇�R2�\��ɰ>3��]�ː5��i2��P�w�
�!��K2���+qԋqg�>�B��r�/����*'�=�&S���M�/0�>U��'��h��q�ῧ����4k�����>��z?l*�f�E�m��7P��[��մ�c$2�2��S���	[��Hj���o[
׸z!j�Q{u5���I��^�
g�ZD��ё���>ֿ�L�*�e���3r����b�|��*og*8�y�j�ʬ�Ջ�Ù
x�iݦу�]�!�p�)�w8,�ڕ�]%�)B��x���#�sW���s���V���fp��T�a*r��6�+w�a]9��V�KӇ���:.��x�]jB�9�}9�4�����Za����qw�S!{G�-i7��q���`��"��Sf��`��-T�(1֛IYM��K!����+C��X,p*ͦ^kv���H�g�	a�ʳ���������]� Ϻ�����f�����I�S���NLgLܤ��>[�������d_�M�����r:7�'���>�~��Hm&C�.�?b�\���]<>ܵ��_��t��XP��ӱIm�*^�t�"���n�U���g&�V�]�.�<Hzu���N��K4L��_��Y^Ό�F���h�C��A٢a+�l��{t/E]`��`�=�5H�jD$��G|$E�!^�8"�z'_n���-8sb����OOKC�4��U��oT�t
<�!�r��kV��VN���t��j�%�_d�s�Rzj��: e�'*,���K�^�Z��+m�` ��[с)�?HJ�9��\�GR �ĸ���+>j=���'B�n��c�߳@���v��}F�0N�������2�Vs�3��L���;�W݅�^U�K\���( ��]�j���b��o�xcP%�u��̭���y��>xq>+w�N�t�yME`8���i��"R�yp^��4l�Xs�p�=�@�M%����=!^{�M<��擞Ʒd!b�ކ����H�[�A<Ͱ3�+��W0�&�L�gs8���w
���:�	�Rlo�
��j>��'W7G{n$��Lo
�}�q�V\2�1
���9�29F�BB+� ~^��� �u��6�T^X�ֽ%t������{1V��K_���h���yJ�n<��ӊ�f�/`���8���H��A�N��O~�#F=���XAk8띛�
ڣ��B��6��mV�BUn�I�l��5�9�Ű�G��6���)]��������'󢿮��7m�Q:�e�s�/D�ZRqpϿ�V�.ԮJf�M�?lQmF��iY���ݢ�^���7�е0���Eܥgj���|��O`�VkEn��r�� 6�t��f#F3�f���y�F��t���Q!M�H����{��JFהH�Sn�6�!������I����������aA�*�w;B�d��zn���cK��j�U�F��b)58�ظ�Pߩ��iN��v�w.�I8���e/$c�5�e�����T�&݅P�������Zb)ߔ~^L�7�*��#��e�0gbSɹ�e�η�M��\�����v\�-������W������徳Vc~��U3!��F�0sY��*l�L�?��ů�j��lvI���+b��\�̠`剏r����/�&���x�z�y��`��>��\�1��I��b�ժ����H2N�����A�����Ѷ��.�bX���od|��{ʅ�e��'NY�aX���4��=����L:��x#Z��%��@�VԘ���e���AK��'�C^q)�P�L(c\iKn��#r~}���h���}h�y\�2��X��#"�HE�Z���W�Jw�kF�Y��ݚt^��C�r��f���XxË��y��ӱ������ g��Q*�|���KvZY:��nJTKӘuZ�%0��/�����_x�_�斫�����|8���-����Ǒ�Q��w��	��ѡ�j��C@�T<ؒ���O[��Z(�*SK��3���:��DCN������F�td?���t&SZ�x6�0\8����B_]E�=Y�vc]�S��!����` ��� `�����6��>��;tF)�4j��_�:9U�x��͐MQ��c���ɳ���;��w��!���Pj������^�"�vZo_�i2���O��ؙ	lPW�2��U 5ե��_K���R0p;�|m��Ǽ=}_��.������N�1z�~�3c�Ds��"Ƅ�����ǵ�$˳���vfrGc;�.duY��w�5m$cZ+����C�Y����]��"PF�<v���w_B�y�В�D���k���M�]�;nS�x���0J����Ë"%���u'�F��+k���jab@�xF"�ӟ-v�����7��}�Q%#�@����t����X�xY��Gӌ �^M���/v+����o�z��D��߮�hy�S7�����# �T0��̨���&���Nc��&���K�̤՟w�@>`=�l!b�46��=H��v�͔��<�K��jh>84��w��
DtL��Υ@�r7��^����_���]�(�DP�	������#�:�82����B ����_�?���G���.!i��<��5/"�{�����Ԫ-v��c����z��H���tK�s�Ӟ��Za՞�Yl��;o��Ǳ��4�V_S91�*o$&�Uv��<q=}+�;T���h��|Ȁ��!Q��rL������+��ռ̽f�r�s�)UǷ.|�*���=�qF�N��>�{B?|�p�j�#Sً�sA}��,;*����XYB��Lf^�D����RO��2Xi���U�n�:ޖ�UMGs�(a&튋ހ�*ļb��\�k'�O@�a�?�jr�G3y�3�����Ʒ|/~���0����pd��[j�����
lg�W=�  E�Kr�Z��kC `�PR��#�4�����cP��}v��M
�����+m���j-��9�VD��%``\^��a�x��6Ǟ�T���ч.��/��WS�����M6�ҋ�ӥ�"@q�����lCZa�u4������uH��U>��s"B9���j�87���QȠ
vp���^_��SPi��H� �LD��x�l5�G��=�r�/���w�OFa�~ᄆG����UA[��b���e��i8<w�d��Ye�:6�W�h86m��H��� ����<�4�`�H:����F5�W���N-$�
ݎ�o�*zd�������5��!	r���a.2L�j8�wbh2�f�6�+���q����L�'�ƢAE�Eވ�1R}+B�IS@��Pt7�+m�~jlˡ�XG��1�D�o�P����P���R�^1��W�t�'��xb��I;��a
�]q�N�(�u	r^p��-3���t���朠��wM/WL�����?��^�zH<�}�V���Ĩ�(��k�v�* �V�"V�F�MnAe�9��L�h�i��)��2>j�
Pv�;��	뻙>f�j��u�*c�Zj���P����H��"z��"C�����S��ϊ�"�3%i���GѪ=a?\�S���� Un�7T����>�9����}T=�4�y�.�sD��d�Vo���\*�����:��X�W$3y��&��\�µ�~�E����T�z	���޸�Ιߏ��q��v1Sӫ�K\���zH�Ͱ��+b���,skN�2a��4k����dY���/����۴�|��H�b;u��'�dic`���w�	MO�M���juG��簈�Ν�l�� �k�-|�<}(#G�����:�td���|xCqv�Ld+ͺ:�Ն3�Vӧ�m�5ڲ�vTP�H��;]����c7���:����d����R���&����'�Ϗ�`I�}���N�h����A�:L��������kZ���@!�} ���n/���$fQQNI��8�/'�'L���"��fo�ǖ�T���*C/����ڙ��Ў?2P:�p<��K����� 1���φw-�A
t|_�0>�ä_��M��>����KdJ`�2iJT� �9G������XI����;�-�.�0�� �1�Y(�b8l@�-7}a����$�>~4K�[��o����'O.0G���H�o?U_Z�4RYɆ�%r��{s�c�jYb��1>f+������g`��0*��0C���A���/�t���\9�1V��c0�7�[o�)=���=��j�S� `K��;��l2����-0���a܌������}�P�c��lX���k��/�k��L(�;~���ˑ��ʇ��f٫V�!ݿb�z)TOW�8,�n�?��sf��r@��-�H*U)?@;�����b�z �K�q�ў-�_Cչ��\t"��2�@ڨ��p������2���ÞG����|�K�6|��Q�*�]�p�{�P�ng����~��Ǵ �+����'&�ص(���#���I�m/Bɜ���o�����,�&��#�F�?&�"F�o��{̏3��j5� ���6{��?]c���t�Ad(STK��1�Y֧���D��>�xo0���j�P���QD��9�3�Ǌ��VX�b��AU��JH�4�u`�ߛ�wǘ�K��pc<?�)Ѭ�T,��c��)�0ZDោ,塭���&��� m9���1e��?ӧ9�����Oį��G+x�,�ڨ��ߦ%�!���A$>QA�! ��"��!øeQ�9����s* b6����n��ۿ�NSϘT�➕�|�׬�Տ�Q�Yф	"��0��$���~���/���,@{�+����c���
w���gu�ׅ=��j%5��N��8e��\����O3�{�(���z�ym����5����ә�̄��d�F���*�7Fғ�ZL���4��������L�ĭŕL��T���!8���d����������vힴ���Gd@H����gH��;y�hA���A�u�ƫ�(��1I׾�T{�Y������)�j��ݴYSiK ��V�/y�5;D�9?���v	���WZe��(��R������*?�[D��y��x�T��'�������h���"��6���렩���h�ؘ��D~dK tAw $N�.A&R�xq�������r�:uSsl��^��[<�)�'�'�X�������&$�6_>y���V�o)�8K�/o R
VgX�(�H��J�f12s](�3on?�7㭖Wn?�V�
k�"�	i�Cv��ŝx@c�[u* WujVU�' � 7��ۅ����rg�76�I�k���e��xa7*�����<�}{���%�܆�����?xx�^�9Keg4v�:��ԏ�v���ǥE<LLwU����R5B�u�W��`�9&��H�'����F�<�T�-��+���Pt\�j2���k	�ş����ك!��?�u�<��t>i�G).���:�c�p��Pa�O d9���(����H��m8�"�'�k�6g��^l��s�ڒ�vg���[��/c�-��;��REhay�t(�S6�m$�A��P��mD�/g�}�Cq_�]?�����e��Q����_�m�F�/M��<�zZ�|_�0��7�{���0��c����}��Qj��48�Р��9��T�_�����M��X3��t���V�c!łRs�vQLZ��!A�>ٲ����9��^N~�O�c*u"5������F�������hx�����ھ�V?�a3Ƨ%wX(I��w� ��2�D�/�%.�{\��7��a��eqY��Q�@g^z�� Z�b���q:gC4�k�a<"j�r�9�nr��0�]�'d[�Q#�ϊ���MxGw������r��N��g�!�����X�Oة
��Τ�ZCգn�p|AKQc�LK��@�u�r�m���,I=T������
|m��Rr�������ؒ�Y��=�aֹ��� =yL7�'d��\L��z��&�Imdī��ŋxy���]��
��q�=y�x��{T�A�Kx�@�{��*߷�67�u��`S�~}����$r���B�/�4��,cm@>D->>M�o�y�b��2b�jG�^�+�.r8���}��W��t?Q�k�;*M�ce8�V`�D��P@���&K�9nb҈a#�aبޗ�Z�L���jJr���o�A��$j>j܇�
�"��Y��Mq6b�*\�8'�4��Jz�������X|8�������U�������Y��1�L��Y"�&zJe��xq�̩	�b∳�W,au"&��-��jw��boUƫ%~?І�*�N�X��)��]�Rq8Ǉ�PӨ�J�%�xp�3�vA��Z�j|�bj�Y�ej��
�;A��@�Ӿˠf�d������.H�:��8��1�;7�C�x�E\����� K���>:��PŚ����e�����[K��v�;N��#<���u��[���4��рR�k_�\�{l��i�8�G@@f cǟ:W5�Ҙ����r�!��A�{fz���7jka�'�cq\>���aJSu�,�g���e{��5� Y�z�	%Y!R�ƚ���G���O 9��r��r?����n� \h]M���aj�;1�1 ���7Nn���o5�C�t�e�oQh0�
��@o���:^sD��nY��×K�����IR�(/@h����g��a� ްot�lj\��w%�wb,�O	��֝4[�I�Ď5
���D�UԔ+���@~��G�q�=K;�JԼR�E�:\.��}�:A<�^S�f��-�0�]^[�o�אDFjBpn�QfN'���$������D��p\��+`qu������^��v�/��vzACV�7z(��s��+"B��,�����V�fͺ�p�*s�v�-�����V�e�v3=��_ކp+�ڬ�mo�����_��cH��H�G_�'�\��fn�=��iR_5p�I����>������+� ���vԙD�][�ֶ����	�.��))��B����׏-.\>2��x�KK9(�ԕ:���J!��C�e5�@�v@��#(\z����¬����Ryǝ}���z6eFqMo�<ގ�g���+az;�Ǯ[�l3-�F�xg5W�a׆߇٥%�xSUĦn�du�_�������,���?Z�0�Z���r���W�2'���1�l�o9zN�j�)�Qv�-Mݞ?�A�'��U�R�ȍ�h�$���0��=��p_��5�N�ڮ-���T�B��Wtۤ	 PV�6�����G�L��H"�R�;��"�yō7 "Y�}G፫!5>.��(�����:��"�L0�^�R���ܥ=�Xb�b����j��No�,T�x򗓽����%K"�;ls�5�T�,�W@XH/�g6��>����;�,�֒+p4��Dɼ9]P�d���
B��z���V4@�(�t�u+���X4�.� �OVBʔ��U����a�ҽ]��.�O�y�Le�k�68��u�5�1���!��v��,��k�~g#�)Ytõ{�i�#3�����j=�u�D�?�XVp7�ac�.��`�*�[��^����nFa��%����.�Ϭ�x-� |���\3��6��ev�;8��"�=�7=��͔�e����������I����4�<f�J�Q�)�%�jt�m�X�n�y�����񰐙��ÐN(�s���L��0H>�/�oǓ�Ԓ��l%�nR^��8�+���WO�6���\h�����QB�Dج0zkRQ��>+����e�	��u��IA�����옆��q�_P0$�T�i����t.��:�!�����*��W&�3��g�̑#�e~gY��6�q+�WO1y_0��2��;ótCk.ZS��r� 9mQfI`}��U�\�>��g-����S�8���<M(g� P#j����q��oZ�ht�J�~������h�T	� �Ԛq?�~��� ��P�`�ԡ$�.e���'c�Үt��0Jӧg����+
,G�K�a1�w��?Z���	l?BH�Û���R��p�=�u��������~Lp�A�cc����{̘}0[�nR���G��(��x�wC����v/4B���FT�q���v��&5�'����e+ᅈU�`�u�HFm�%��_��CM��
҄S>Ǫwރ�<�B~��52�]v��K����ߓw�����(����\�I6�2�ñ.f1��t,Xv{G��@�8%̯�x�.i���;����ؼ6'�aY������s0b�X�QQ1ekpS�]8�6vP3�>����:ƅV�ǵ�O����|t�ӘW1�p�w��*��i����8,�K,���0��/��g=GeVHU_��	*v:)���a��6��w*`�Ұ!�;lV4�ņ^#��!7ХI��B>�T���r^�%67d}��=�=��Y�ZH�:�s�B;�玭y�}ƌ��T��r������f=(����i	2�)yrDk���Z<g؏��)����B�^�xt�7%%!�W_�5ս�D�s��,�]��F�Qxl�����M6y`��n׈�Dg`$�]7���}Y��%z��´<F!����l��I�
�S��ܙ���~���܁���W�J�y�������1�'����wE�5,3i%� �Z�2�*�w�a��?���~%~!/�)��ȊѪ5��F��S�Gl��3�}�&�ׅrI/��;���4���yI^vGd�85�e�T��%�a�vJ:D�/t1�a�;eTL��>�*�5;^pB�)�������������fX��K��|�v7w}(·K�jQ�ILB�/��A��%���;��BUc�I��j�kS�µ
H.�4i�@�)�0��6�������#���x�����ѽ.,�x�B1��Rk>��p�J�\�jq���/��z�\$l_��Ҵ�X,��y|���R>�������b8� =�i� D�w�c�'�.2>1^�;��nO�%,i���d;��=��4y0T��2ݥGa�[�ɨU;Ї,����b�S�'q�ӭBJ���%e������)�T�&�����,�)�L��W"]vr���FJ��x������_j�l����+<���}
\�
�8�����b]G�����4@#v��'Wզ�S<���;[��?� ^���-q�Eۣ- ����@Y��+�:�M�)�~���~�� ��kE
1�x;;C��2�h������i���X*^Ǖy��T��@#�}��U����].K�}I�u5O��h�0|�I�Ō`��]�j�{'��K�6��.�������@�p}��K�}�����p�wq6(v�AWR�!�@�{�zZ�>��󛏱�6�������@$CΖ��w�h"�O{`d"'��FY����ߠ��������߫|�N�I -GX5�A�^q	J�_A�J�^�H�ՑRP�����s� 4q�;��c���N[�{+љ"s*jA����CllʃF%�>��5�=���)o*�Ϡnq��x�����τ$Tz�9uBA�����;�q������XYX�g�O�O�[LП��CEg��[�%��0[ ��r�߂#S���	~�@�E����4�j�ۡm��I�G��b%v�H��ཛ�Y:���na�(�	'F:��)�%y�2���kzv h��XwE��
/�{���@�( S:�������m�"u/�GKI�q�d�N§Y8�n��lm�3�e���S�  w�_X0��H�)�v�B�*��t���v]3�B�h[����!�Ct�M�G|G��4AC�7�I	e���}����n�4d�2��j���ѳ=�K}O�J%g�X�71{��}~˦��_�i����"Ţz�L==���H_f[pE���|D�*�Sl�������)\������q`���s�ƪ���;G��HI�'Cf�dεM��4��F���������X3kk��z<J&4�q��!i�UyjX|oB�c%2�W�M��-^2&m��s~��^���m�2��a�p�U3F˱9%Z�l�]��e�N�Ec*�߾PRl��y�m��	���S��P�(+1ݞ�jK?-^?CK�R��3����\/Q퍲��2}K���k^.��C����r��KU\�����-RV�Xm��q�i�^՗/��yE=/�Y��F~+���'l�/_��"��$�' ȹ�1�w����#H�B�V�s�V�L�;�� 	
�b���IVh��׿ߋec�a�����3���s����z�dBj��G��M-��w�j� g_�k��/�����,�sk-ҤN��E>r��~	�ݼ^��!j��"Qf�n$���j�>X��xuF�f���X�W�_��X���ct�.2t��U�Gĭ������S*w�S�9�ϛ�v|��Yfx"����?$#~H���=�lΓgX8x_����L����S�P�eo6�M� ��<�W���������b.3$8/]"�֣5 m�	`F�0�+t��O���cӭ���|$�z��a�����Q&+�4o���S���@���E�m��9�#N,���
[!u��Dzj7��7;�l���ߋ�<��H9�?dx	T��Zŗ��� �Yt��S?Z@��R�9WĘ5*'��`� 'm��+�,�2�+W��e��7'J�5U����;�J� :~�5tm_a�E;\M�&
��וk�|t;��|'?�>���yl��ƍVGl����f����)Q����z�!C��F��W^gJ��G/���W^� }o�E.q���M��dD��98��rϽ�%����9�����q
�a�ty!ב,OAh[��0 ��@�<ӣ��7�(= ����a�,X��J�XQ��\]h� 2y:�
	SjO�U�puX8��2��`��G~� o�8媫 ���T���A���C/�l�x;!��Ә.�R���l 2���iA`-ˁ���3"d7�uLȱ�pB8�����K�Ɓ7�5���~f����I{�P��r�0��
���ꉋ=��{���ͶFN�9͎}���F-}|�A'5�֊��V�=(��1�!��vԐ�8���tMt��us���#��;��rT�t��e�
;r�H
��޹�%2E �ú��h����\G\� �jš�3n�K�)�	�@�Ӻ?��7GZ�KE��{�KG�� ���M�ʞ�{v"�h�yOR%BDB�4�.�����ޟ����U����xo�ǞW�*à§�ӭ��׀��6�[PW�&x�5{���4�2�we0�-_�5,j$��P_��gd>%�8y��B��y0&�R�O3�~��Н-q���}ܬo���^,O�D���(�Wh
�>g��]Z`���#����H��T�>k:���ً�<N7����ΰ}:pE���?&n�1�����S����s��,� �%���S��)��،��|O��5�w��^r��Oi��"��d��Fiʨv�_��o�8]ι�C�gŴk;��k���r�rU��5���2 ��a�q���襉-�@�� /��_V�e����d!��H�DOl��T珻��z�(S'�Æ'�IZ����Tz���D��Ū�+��nM+W!奟c�7X�!�V[Ɗ�\�h�ް�M66�s��{g��Cq�L`���I�qSf�Sx|�`&)_�0��#�����E�g��,ّ��|/�h��V~A�*�$u�]�|���x��k�A`��U��l�?��q�ѕE��w%|�NϸԇH�!z����I���y�p3�#,�e�.gz�m�Cԙ3$��,�SNJ v}��ր����gЧ�L���f��D���Ҷ���jgN�,U+�s�+�AU(�m�ީ+�\�G �ْc�/y��T���*c��g2�%fl,¸:�s�M�8[Gd$ɵ���W����J�N�&���_�m�r�����@3�8����(s�!q�\q�)�n[lM���~S`���̅�#EA��=�k쿵nvGpk���*#"Ȣ��d���^�.eB
����|#k����v��߲Q ���H纛���ʖԡŪ��&�=͗�pW[/E9��&�,(PS��{uKjnߝ=>�Xwǿol����"��;ZM>q( ��e�`�:]�/�
�ڎy7��M0�;-24�׸��\�M�B��"!
�nG�:<*t.����XaS����};��S���2��#�@n�^�廡���S>}sEdp�������gx/ 8���A�Xi���Bۯs��mg�m���a���J��7��4Ϗ���U�}\؛.�9Smc��L�4r�m��A�Z2�}P04��	`�6�X���sũ�tR�}��'��U��NN`�_��pKe:^o�����p�7A��	��;�N��$-o�5�X*��l8%��66��m��֬�L��<
���'h�2o@��.Lt�]�#�ll�vڦ~�g�����S���m���f5i�Vr��1����U����
��1�.͕7�������qӧ6Ѿ���cHX�,����[2ī��(�2�t��&!�e� -��!?C?�gi�$��"�+#� 8�:L c��w8�q�Ӌ$�n����h�*",������w�\	�Ja|���V?�!h�����'�Wh��N���뾭����	�0�vBFC���#K��3�����}MO_�ƆhH	 �����k�32J�QΕ�۪_��$�o$����W]f��E&
��Xc������T@�(R��0�D�11}7~�� ����;�Q����g�u)��[��9��o�D��mQ�ܪhn�pZ����'���S6lW�T���@�E�9�������
.��D\
�&�c��!?H�hp�G�԰�"�O��t�u|9N���3�����zJ�ïrI���k�����~�v�#	=�i쐈��c%�z/�5�6��--
�3����ԛ펚��1s#x����>�l'Y��s��V^�����g2>� ����������G�̔a��;]/��fZ�(q���T���um�8��P�K"�ׅl�,I$T��Jv�L�T�E^�.,L�`�Kg���)z?c�CG�0�6�:��+
����_��z=Lʔ{-�.fX�#�\��n���ڝ�rj��;X�%��g�	��զ����*�|f�br2}:U����T��X�^,����cr�}���a�-���������Wi�� w�C�i�(�<��%�*`oPΑ����U�®��
E5�^�Wuq�9��*�I��y�;n��ܮ��J�zY&��y�J��[{����H�IOw�az��aF�NWJ�}�'��*]�/kx��*s�~-U+c[��t�I�jB{�7�As���,��R��l7�c���|�ڂ�tZ��Ӣ�������X�<�B�a�Ì?���p;����6j �&Ds�ta�d����l�}�R\�D�U���Ǫ�J��Fݠ����6��x�|��>K�I=��ʔ�����.XvC����'g>qk'�1���,k7ܺ� �a�S���{{�U+�Ht��"�*�ch��y�xU��˲��N.����vD�{����^�'@}@("q�i���'7� ��Ai�ut�1��]�n2]3�l|}���S��a�ץ����"U�L���L���.R�#[Q���20����:G��$]���ֈ$B�.V��`��$�{���7a�Т!,��}�4��Tc,������\Ah�PK5�8��;�%�U�h͊���U���fFjX�M�� ��'t�����W���o�k��dT����D�2)���m,�D#�-X( ,�z&�EAҺ#�:�D����!�AS�9Utr�_{�# z����G>�)'�Z+u	���̏�T��Hy{���# �y��6�ւL���)��X�u�1AX�*�[Q5O��L��(�.i�Hpe|S~4q��_a��K��	��n������&�V?�+XM�3g�\h7��6W�&�l#�0���bpV~��������4���$�f* #,j`��kZ����f4�;Bk�vP��oK�װ��Ϣx�f}R�!�K��*��?BAdE�
1u���W���8ض��ݙ������+�`�_�\���R!	�`&L�`y��8"�ʾ&'���^l4�QzƝy�M0�Q���uF~�K�=,��z������3�\辰�݂��ar�e#L�eV�W
��(v�.�]T���\i�ۃxmƘ�9X�1��m �͏2fxޗ���q�]��0 U�.�������s;� ���'�('gŠ��{�|�9��^	'��g�FO>hcU�o%H83��~�U�#��f8gA�*�gG���FC֪P��T{�T'A�M�C�!0�����4NJ\)�w�DG�����2�|��
��+ E:��{T����-��=)x��AC���4K��{�o�mODF��;�Cۡaɨ�f3�h'4^z�jMqH��s4� os���ԋ1{)����~�<ߺ��b�T�e�U�ry�|}(���n�� ��G�.��=m`ݣ�1��)�+<�L���kd~ ~{vl�?5�,��#:�Պ���J����f@�S �b蚓�U�Q��0_���D�8"����?X���9���{�"��LPOx3b��Ha|QfP(��m0���Nr(�WB��-1V�Ɏ_a���Q��֪	�,�s�ו�ғ?j7�z��ڪ��wm��L�ɹ��U�FQgӽ�_�or�'S��m�[^kx����d#��4�~�օ���^�+�����K^^�I$#��	Brs4��_~��cֿ�Z1J���-�ί���C�0�D�������(��$����MF����5�'�����R\ib��  ���[�b��~)9��Z�|�7B�H�-~���B�k>a�Z�c�3#4����%����-t�ԩ�I�aS�[����͎/ ����r���}X`k-�����1N�Cc��~���7ȶ�]���}q5�	*��W=8��l��o[׸�=J�Y:�4�T� 31򛱋�h�!�K1��p�z�zZ�R6�?�.��Xx��L���{��I����
�y�C�J�4>�t�ު��=�&�����/�%W��I1;;��v����g�X���ij�~��G<�sĈS�Y2�^�J�ZȒ}�O	0�R���Z�vD}������
�yo�UĜy�M�f�ϳQ �#o��x��#�`����m,���}���``v�t%[7�|c���*���-9,���2͒�{��؈`s�Jv�(w���k�4�L�\�=	�>BJ��kuRz�v��^s�?'i�?�*�tR鳆.�B�r���qP�[Q�j>9��)x �+�1���ԽB&�� ^2S+���ر��'L�-��H%T���v�?qC}5�����V�y7fI#h�9u�F����I����M���<�qd�N#�}�$3�,����.��b��&�_E)�$�o�M2����R͸q�0e���7���u�����OL�.̈́�P8��	o���X#�H "�E�xk{����i�������/
7�X�z!+A�p/��x�_��9�
/�C��5�a۰���x0�b���c�?{�?YW��T)��P�r�l-㱲:�xkt�_EW�O�"�hc��+��3�4U�[V�7%��N�o��헰P?�2��F#ѥ 8i4�c�[~We�Z��w����~{���N��.q����|&}:=GH��ǯ���^c��	�y�4�'ŰO֌�CW�o��R��I{��x�nY�o>
�����=����vbV�����"� ؏���V�T���q�=��:��OU0�������z�<_����@��0��u��￣B��8M��<O�?t��X�L���S�&�O�N
#�I��3y����������\W�?�
2\(x��1o��y��is�Q�P�V�E5���pZ@�� 2����\�E�:e�$�aBX�-�ϫ8<|�<'	�M>c�g�\��M�[�T�H��;�6�,3$P�I�Β���zfEfo;�lZ�"�u��(kI��Jd��D������ a6�i���D^����H���pe�3�[%�J�.��g��dIW�^K�s�/F#	3�.���B�"����J[$�e7�g��h���eғ�D�2W�<-b�'�e̵�60(A��꠵��b�65����-J��:܅�a�:_�zVm��e���DPp�t�ɫ心q�Fa�Wh2�N�$�:"��A�c��� ���]U��-DKTJIoG�n���U̲����7.���V7]L�h3��l%����ZDB����w�g*��8^�.rh3�h��x���䆊]��={L6Y/6 ��S.-��}T�$9������A���F��`���A�5�����Wa���d�'�����9��
�e����\�>\D�%x�#�-�xÑ|�͈�I�q��U�\��
h&`Ȑ����h��Gå��SN�9+���S�����{9i/wŀ���(�?��\�����n�YKpγ�?�8xz�a��8��r>.�=�3�44L1fH���U����f�M��o��9��3���L6��?�Ԉ�X{�Sd-���	��E�h_ώUˁ��h�>�֬Ǣ�X|�-��*ˢ�5�� c<�ʍ��� E5j�$��2�X����"�[hL����w� #!��/'X���+�[�F��I����RƱ)gr�rrv�ǕM_;ˈ(@�n�-��`��]��������������ǰ110S\��2���������������&3��R��������Fӧ���p�G`Z9s���B���L N� L�۞ɏ�Z�o�-v�2P�1�k����N��zk܈�(Ћ0R�9��\���lDD>K�)�kH�.�'0թ���Lʃ<��Vb� T� ��m���j/S�>��^i����.3pҼl$u���Z����3>�n�1k�>���p��I�C:��D}��I N��sȾ�9V"�16�R�9br�hY�EYt��!�JRkѭ[ݕ��B9� و֥p/�˒�!���o��x/�81Yl��qI9?[f�-5:��U5f��[i�T���K���yu�Z�s�P�7+њ2���ga��D���vQ��fv��LL�
�I�5�D{߹�a�EG���Q�?��6�`h����y�[�l��^�I�!�=��rv���0���Qv�+Ǳ��1D�̑ٞƬU�y�u��mg��8�9W>����[5 4v���w�r��q����--��M�I��x�-�6���ϔ0\�8��8��J��d��)�/-k�������=Q?�J�-h�@��]"p����p�Rv!>}c�Q0��mv"�E�-p< wV�[�h�����Gr$r3��Rqڋ�kѹ�3�9:@�biwc�!�͊S�g�7�� [
��);FT�=5����ۗ^�aݩ�ܪ�
��h��B��u#n��M�E�H����'O����UK"�{��dkI����u�w�qh�uᑿDaZ�&1F(���e`m�����r�`h�D�"�J��T�+S��D��yg���bɻy��;N��j��`o�j\�tR�a�C�����׏��eמ�����r��bM�Ҋ�N���(	�x���ߚ�9�q�ɻ���TU��½=�Ҩ3��>��ȸ܋��׸�R��P�⩇M���|ibD��"9��"	8RwQrĺ���@���S�5p�/S���y�%��}�ߊUɆ�Mă��+��2?0�҅\�]_�ݠ��1��"�d�#�C��(�ܩ;4�3b�[�*����D��b�(��-y��%)���°][���w�
P��dg-�8|ҭ)�B*;)�q��8�q����j���A}%+��1M�����O���Y�$�x��O��c��=v�Wp�xu�F[�s��+�[a���V7��,Q	��Y%�[���:��Yd��D�\���C3Φ��4��޾)F?�7��N�a�Y�P��[��I �v۷]�D�$#]���|���z�\��������٥�q��u�لFi�9�7qR��Ԣ�;���ͮ���	�����Z��I�ڎ�����̳�I+��Oe�M���e��L�sг-��$�U���@�׋�I�.���pS�����F�� �o���	_?}����)M�3�7��̜�]�;O�A���ȉ�ˆ;��ʡJ)��]z���3C��b���E�_iu�*��N.��uwn���4qS���T�Ň�+�/�rc�͊�zP
ē2I|`�rP�����'�^=���7��I�y��u{�Ws��A�R.�O�t�ǉ?����O�o���YsN��i�(7��CB*㜮��tR�t��'A~I�d�vhYC�O�f[�x�'HO�Om5�����\Ҟ�,
R?�:]��P��Џ��+�~\�c��C���ܔ�QO����k_IoSz��6pl�8��K�8��b���2��%J�1�S���������]�w�:,�?˸[�ǽYNl�����B�B$�.4�ł��{l�fr|�/!��P8���vRQǪ0�	'�@�����W����}��
�Ŝz�C�5�_@�Zޤڡ�OS,��5#��!o<�U�) $���lY4X�%���}l ��79cco�U-�ϳ9�Wɸ�йN�u����!�K#�7��<�~W��i�!a<��}ߎo����&�������1j�����̖+�4	������ߣ�%���>t�gK-�`K��K�FK�p�n���>��x0��ȫ����Ϭ=��;2��%�n�P.��+Zo�~��p�<��5S><��iQ}�O�ڮ
���&�A)�/�����p��9І��s���vC��{Vt�P�����Kڼy4Y�gl�"�omϦ�o�;��I	u��KD߭ ��X�W�� G�蜛��4S8 �N��ŀ��D��(Qc�;�A�x Q�[�n�m���n��8��`��h�A�z/E��3����j>����A)��)�p�3U�"��Fl�����{vfa��J\w�-���C0}n�m�w&�h��N�p�J=���OBC���<�=1�6�zUC{�~Gԣ�@��N��2B�P0az�8��Z�.Q#e�5��X�}��� ���B�u$*KP�й�A�z�������-άf9[Ko{'�>��� (�Qz��.F�v~�i����E��*,����g�rX.�x,�x�����C�G5,����^F�]�8hM��k���h�w|�2	��Z[����̵L��V���e}�Vӽ���k���kT���k]�4�����渠��ˌ�	�-�r�d����6�q5���n��N���m5uSk�텬fy�3Y������޶C�_��	�mp�=��2_�ίD�7��j��HgwJ�9�T���;��ԓ1�r��,Ȣ�*ʃ�2�",4��\^zͻ�0���¤C��\Y�'Âg�-��xpK�tB���Ѵ��L���n]]����qj���F}��%�c�j��`-f1 ���V���C4��:$@N�E���8����M�7����Q��7�PҊ3d��ޜ�]H���{O���Ȗl,o޲�C���[��J����W����,?YYƄ�9fUy!���l�K��qfH�T R�A��դP�0��i�{,G91f'^J��c4����]�����u��enA:�xo?���N��Ta�Œ��<|��l��_�>4��u�Zi� `c��[��!~���0�дFi�]���L����Nz[���%���b�`�����ps�s$��Ob8��v;՛O����?=a�"��}ԥ�7�a�@A�L��pl\�
���)KЩi��vf0~!tqn��a�ɬ�����9g�\�*��V�d��vAm�@Z�wfFF�^[W
[��aj�m?}�΄�v�F� (�b�ct]���]��y��k�]}�:d#R����ys�ښ!�X/��S�I-Nr�(�k�%��xQ
D��Đ.n�,r+�Kt¹YMiX���k	���R�ܣ����1�w��K����A�2@��
�P;��@D;���2��a�|`w|�_ARx����zY-��	�;RYg���� ��U��;\�������5��^�Ź�g��kS�`l]яEq��7A�_=�by�'80k�q4��E5�Vi�R7c~�