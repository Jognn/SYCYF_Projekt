��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&��n?��1ů��> K�-� �&�T�Ek/ֆ�\�놭5�DꢘP���+L+X�4��J��#�0�8���������l��jT��+�(���������6�MC!D�;�m�퓊D@v_p��䙋ⲝ��C_�6�Ռ��#�� ���	RD�4D��畓7���vn�H���0���fX����4 �CS�C`{��;�L����li��� y+����FD�p"��]���y��R��K�({� .؜M�������	^5���ɋ��&���&�@*���
e�� �t+���
_6��O<��7f�M��u���m(MrN����z�jL���@T`��M3��c�uQ�Y���%�dD���,�~^���y@Ga��(����C����	��G�86�S$��ɳT�ز8���:r��/y�[ݦڍ#A�����i�&<nU��<[5)�Z�-Ĭv���0t���d���"_���:�'-��d��*��q����_d�y�N-��~";#��������Y��؆���	6ZJnԷW��έ$Y�K�?�4���L�w�Wmiɶ��Y�?jx#*�i���F�m�E����O6T>]i�_�9;�!(��kH7�OS��_��[-M�((��lO�s�$�g�x7`��ZV�E���F��,9�j	@���]}<�ahb5~ãdl&I^�	v����-�@�@���	��!��d��`j[Q��� r��;f�i�.�m+UH7��/OV��c��������l��i��M��*'��?���G� SK�M��H?�7�|��}qz)(Mx�(��CY�5դFfa������Z�v¤[��n�y$a��̷@�0��#���^F�Q�*��H� 0�L��4�)͉Wb�e������ܴ��N.��M�h�('�o�ҩ�@���~�@��-�}�q�R'w��1�*�b6��L�C��5��\	Kg�eM_�����4*xkw�+h����R7&-�X��p��?P�ה7/c�2}'?6�<i�xԩQ�?�t��#�H�M��|�7=�(�y�+��ݤK����t��ߋzf�͊��swT���ѧ���e�c��L��C�����<���+P���̤{���0�)��:��'�	����&υ 
VA�(���l���q큾郣c�N&;�F���Se2(4j{L�-B�݉�4��!����E��ْZ�;��gW�#X#y��N_�b&'Q��ZA:?ק�*��|��Am�Y������5EH�N��ƾ('�K�4MzP�w_����F�]+����Dh:�D����y��Β^e�zf��*3дW��a�-�����o}��F�@u���_x�3'Z8Z��Ba7J]�<��{g��H>�U�Ҁe��X�]G��� G��/Z�ZT���l��C
�@��g�H1e$�9�v�|�ӭg/��\q�Y���R��!o���ʜx����̶��7��:��S̈́k��$G3�f�7�I��X���J��l��ۃu�W�sM��F�ό[�3}�߄��U���za������gA~��Q`�\��o7(n�D3�_ޚܛX��Vy�A����f���@�8e�t���S94P����Y����1�{�*��`�
|�����3=�?�]փ�$.8mQ�Q*��Ǘ�-�z�ɀ��Ya�v\]�%��������_���ҔU:e���>��x*O�.�\A�g�ވ�I_TvkLU��qi條辭��F�f��ƛ�A��q���G����B��`A�eWM�7���@=�	n� ��	c7gJ�;�(f��@�+%�e.�`Y2����,���vb�\�y�F�k�U����g�u��C���
�P�]v��6a���m¹��%��z�ːB�n#�ӿß)��é;�ş}z�J*��$:�������L�ë^ P"
�Kl���z���T����ˌp��-���Kz��׷�Tc�X���-̶�/^�T�Ej@@~1O|6�#�g�� Yr���4xޒ��v���6y�z�N�n���l�'��о'�T
)3Oi��V��4#�6�}�s�|R����=*���g�aѾ�L�拏�{E�~��B�Cɓ�$�s�y2 �����Ĉ;���mۼ������ �<�@��;�3���Y|J��/��C����q)6!j�x��{�/׬��3������h�w�UD�?I5J0Q���䬫l�H����
8b5Bn��(u� ��?`���>t�K,�H~�Ɖ��,#�Abc��V����Tq� �9� ��i�5�ƪ��s�)�\3�#o����G)V�k�k��wv׵����}Eq�S�� M rn؃���_�I����`3mHg���"�`�d���|�g����pw�ә��9���i� c¼��_Ra�)�1-�`A�[���E����r�<���~
#N�|�b.\:;�D��}�Pt��{L�B��#���%��!����5n�Y��m�p��_JY���� $j�p<l����6�^i�#�*�F	6���*X���5׺X�y�]	�#!~!E�\��zz]��f'y�
x�Ύ-"I����L`5.�� u�1P˔��!���k)��M�K�W�qM� �=t�/���76P�|Z�I�������[��)x�M�<�\�c���-7X%�V���+5���WU�I��ʈG]�҉��FwVъLU7>�'���>�c�� WvE&ò��l���P�p���?<;��W��u���4�d���NͮTI8�
P�+���C1�+>}��^���b�X�Fs-1T�)I���*�%���_�9����c*������E��u�}]���@�,~W��u����'6� L0�S�RC�r3�)E�U��Q�rDe�-r��A�ZπrԂ�t