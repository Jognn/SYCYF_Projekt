��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&��n?��1ů��> K�-� �&�T�Ek/ֆ�\�놭5�DꢘP���+L+X�4��J��#�0�8���������l��jT��+�(���������6�MC!D�;�m�퓊D@v_p��䙋ⲝ��C_�6�Ռ��#�� ���	RD�4D��畓7���vn�H���0���fX����4 �CS�C`{��;�L����li��� y+����FD�p"��]���y��R��K�({� .؜M�������	^5���ɋ��&���&�@*���
e�� �t+���
_6��O<��7f�M��u���m(MrN����z�jL���@T`��M3��c�uQ�Y���%�dD���,�~^���y@Ga��(����C����	��G�86�S$��ɳT�ز8���:r��/y�[ݦڍ#A�����i�&<nU��<[5)�Z�-Ĭv���0t���d���"_���:�'-��d��*��q����_d�y�N-��~";#��������Y��؆���	6ZJnԷW��έ$Y�K�?�4���L�w�Wmiɶ��Y�?jx#*�i���F�m�E����O6T>]i�_�9;�!(��kH7�OS��_��[-M�((��lO�s�$�g�x7`��ZV�E���F��,9�j	@���]}<�ahb5~ãdl&I^�	v����-�@�@���	��!��d��`j[Q��� r��;f�i�.�m+UH7��/OV��c��������l��i��M��*'��?���G� SK�M��H?�מqT'J,!A�h���'� D��G�T�>��tw�ܻ��l.pRu\7�V-�T�V���CS@�ewf���H�*�cwl�H��ϋ��#�`IY�k����_��U�A#���z\�yz�~�cٽ�bl����S�&+s#�V��%��ӧ'A�N��qT�7a�t��$d��]sH8�G�?����i��i6�ˋKl<�O/���	w�C��:�D��]�l9�ތ�G6���Ccyg9m��<%���o�m:|0�\)!�)�2�*�y�e�M��%����� w�Y�.���,���E�ٗ��N�*��O�zP�i8:³��v�\ݏ*�P�?���`�l��F-U=7�g���w��ȩ��$���"5��!������{Kh��������k�$V,[No�"a�K��H��c&W���Xu3ѳ����i�uI(of���p4<t�Xzf��4p-h��,����<��W%P�)�������c�%w]������"� �ۭ��9�[�Z_���K���N��� �{����Z�@���k}]�s�yR��݋}�k���/���7�&�<�V�0��dG�z}af��5#8��N1�M ��Tl}JĖ�B�	�}E�}�A�	K����D'�R�g��=	������+a������%s,^m�����Ԝ>�m�����?��/ ��#]>؊uN�\���0}�ڇ�T���cj~9�I/g�~0��1���'`p�4��w�:�)�W�M�^�p�r8�^�XO�>j�̫h��BZ�T:�x��z����p<xͿ`����u%�����HM��@\�(��'��b�#d�O��b�i� �SY�L�Z
�=,��H�G�tu�>��^<�Hv��o�z�@�(&\����F��Fq� s�SW�Gv��/������bE���9b�g3D
�'��}d��s�3�KZ�+J��#ӎ���<0}����@A�k%߽����ș39���G�Zx�D�\i�i��6gP���80Βw4S����ZP{N�o��Lv*up1N���[�o)}�"�p-�C�	�,i����iq�z�\3�	�zȧP�Ӝ�n�����;��yq�W�M��BAjT��|8��{]�NeċV�h����!s>�@���Щ���໨=S���p��<o��ʔ���`*�Z�瓡�N�ԯ�g�mo�E��oMb�qc�}��b�+�]|&�\N=�%p�	���"��ۮzմ��M7b�`1r�:J�߰o���y�1��yϞ� һ�����ņQzV.^�ֹ���j�s�qZF�� ��{�`����OB!p��zh���M�:�fH|���01oX����[ԉ�֋���S� �����G��^<�R�_q�zlJ��*=�xٍ%܊�*������V���&� B�Q�M�2w~�.O�*S��`ns�ǖ������{2Mb��0�K�8�o�)�{85�P�.,��~���w��؝^�P������o����h�.�/���%��`��AP��X�����������D�����i�J���LɠQ��e��4)S�i�{_��vXI�Ĭ�_0�)�c�&V�?_���8��xz�	��V��<l�� ����v��b	�5j��w����A��b�V�he�#L�O(l�M�ˢ�`��r��fv~h�V���B�}���u͎'�~(uC�
�1��e�0��<ɉ4pX�h2�7�C�t�6�y?�K]~��fꂚ �z�%PϞͭXy�(�Mw1��y�)5�94���5g2v)��4��ܟ���'�G8�E^�6��#��3�[@�IOm�í��,���fm��Ij����]�8�t���C�9���4`�a|��������MMz�CJ�-D��Y������?>f�a���3��S�̾���m��F7o}U�+�'�Yv�s20�\�=��+y޸;��i����:N�(�ǿ%�z�� �Q;�a�|ք�Y����H>$�C
9�%{"�q���u/G|#�G[�7�;�a��E��d�C�ۧ�A�����K�n�5�1�6J���o��)>Jt�2>���������6}YcTNxg�ǃ���Z��Y# E��g�����E�*�c*^�Je}��N3n��Q8��i�.��N�]�Zw^S���_0����2��o�4���c�^,���ё��.;�@II8߅g��R��Y����ɨ;�CZQ!�jd�ܒ�x�%���"OLg�M,O7��j#9?m�%ʻ��'��Ck���s�,Dh�n�{�M�.�B�S�vv=T������lfY&b��D���~��ú�F����I�C��5c��Q�ļV�D>�r_-J��ga(��Z�B�QGA�B���ʓ�l~�OɅf�w�����so���x��$]�z����z��h4E*(찋*�e � mђV����(���W2�B铫*��σ�tE{ZV$W����M�a��9�����__�kћ��Ϊ�3g��ɡ�1����nûd���o����؜�f+�����v��uJ�>PC��v~���h�C3��
ۚZ��	�z�Vl�w˲���P��6Ÿ�����J������%jb�(��8f�s�Ϗ�͋��Ys�
x�A���L|���/��tb����a_
�/��TP�v��K�nyl)L����ߚ�:�;�+��ȗ�O�^��<����� hߎ=�F]�,�Ъ G0����ȹ�Pn@@ld��Jj:_���ۏ{Z��@+�F�D�N�x�io�df�[/��g��^��.����r��������s�.�|)�b�e��6#ok�2a�YD=��s�a0P�\�:�Z,h�>�= �j�z���2�h��r�):X0�tD����0�`��X��i�	���H��x"P�(c�~~O�[��i����C�ޡ�_1�l��P�:����\�����_M����ɗ\㕯&��k�&�Kin-�!�{ VJ��3����gP�J���4V���Ϸ�:��=����qϚZ�<"��Lѻ�`�p%r���~q���ڮ� �>X�6�������y���w����^"h\�8F���Դ�� �z7�%<�(�b;G���mð�X�И�o���/[*���]��DN� :��#�)�θ�����G��l}��i�tR���L��h:� ����ml�,�����C�����J��9�%��&f%)���`Y�0C�+��i�~F���s��F�׾�{�qң�qO��H?{�u��i:�ڮ����/I����d��x��-8�yq�%k�y�Ig)��]��8"s�ד����������!`)a���_��gy���)�vn���!\��� ;�<bӁy[dڒS������QO�N�~��Նt��F�M��&��o��gG�W����˘�Ԥ���h��]��r�&	���~��<p�p�\ɺ)�}�G�ӊ��\��y!��8~A��W� `���i8:�dWD�zT����������!�śd�Xd$TMd�E�~0���ZQ>��	���f���p������Dr��@�k�b�egR�Sk�f�)mwD��y�Q���I�|d8k�|I�2���p�T(x.Wt��J�_�U�t�1��莚@0�:�ۢ��GUFN�����>(�OQ5aduv�(ٷ�z� ��S:�Ӥ�!���R�r��y�񹙓���~��� F������;j����Ad��Lk	��V�L�!��~#7��}��+����DLMhr�[�H3��M�Ԏ�T\����~�F� {t�'86Aa��Ĥ]f�
���W��N%	� �D�\*=O�u����W�=�ߋ��56I�e�d���U��Fþ1�����ͧ
���h�?��^�>��o�W�[��_b`� J�=����fAsK	�?x��q��]&FaSaL �y����=�����q®����Q�V.|O��օ�]�@S��r����qQb�l-&���Wq	����O�����ÛO�� _i��g�F����[�F�h��)�˽�.�Eu�'�r?�Unl��EV	���<de��}xPf�������n����S��i�u� @�L���]��s&��弙�ׂ�P���3�>�s+���וߖ��3���r[�P���hC'lx�t��g.��L|�9���k��� ��sǁHjkO��"$e�0xQ^���l�p�=�^�gv�gM� �����]�S�t�@~��k��J�G�d�S�cnx��=�?���f�4�T:�V�N��OG+��eƣu�b���U۞/��e'x���Ep%cT���mжu�)��0�RagLJ�SH&�nGL9�njP�!��v�[�?~8�Zl�Q�fs���/ج��&oD(�b�'J����ƴ?���r�8`M���0���é�,n_,jn�[8����K$�H���_ZǙ�^�:ƷI%�Uu��{f��|�B|E��Rh:g����� =6Q�����UO�;%y%'+ΤZ�4�
۞�﹠������c�9/�ȜOD�o�(�����6m�U�����o����������z>}d
��D�V1�9�%.8�5���$[u�)�)U3���k��oqJ�ݱ�1Ƈٺ��Y	�3���ߧOe;��Ę{�e�}��9��>&����2N+	f�#*Z�I�D |f�d����B�ý�H��`�e����Z�x�-��ϧvw�����~%�=��#�tκ�'�i.	�%��P�c��>D�\>{8rT#�� ��^o��Ji�õ�8.�aq�x�0i���V��wx��˘�{r}INT<��p��������ªZ	R��3�|�0xjL�'�ќ���w|~Uu.���+��7��1�����V�F0�.o-�d�K>�*Fs�����Tp�Ń> ZJc����Y瘎-�v��L��g�Hi�`�]�Y�J?Q�2�E*���4׸N�[.X7%���ԍE�H(��"�׳�|�r�_�W�}X��ֆ2�G7%�UFJ��Rǒ:E���-HU��:�3��CT{p&�.�F���X��(�W������D�N�!,�a\{��e�vZߨ�5ە���)>E ����$/޸Mmt�c)�f/$�IA������Wa.N��(ħU_%ϳyt�0Y���+��� �~�%͜�X��,4{��)���|.�Y�Eq�/�9[��c��qW���l��3�
�p��ef�3A�\Μ�B��p�1b��C~��lp��48�%��/�����J�����U���_ �A̺�J�����x�Ղ8/���(h"��7/rSLX�ث?b����E��C�H��x�׵�+�J���-���zV�{G��
�B!]���W�z&L�%���Q#1��D
@x
�$�sP)HK�-68��-�>��0Y� ��M�6jjE_Y�XOZ�D�|�.�|���b��k�K��.7�f�0:EB��k1z�M\Z<jz�F(3���л��)���V��!p��N~�L|7��š闝`��=:�u��+Y��̠F�Q�C��5�8J��	s�/��cu�@*hf��A�wN�ζ���:�@��rB�'K��p��5R��âD!�����:y�`��X�XT[�� $���b�{��`��#5` �L��Q8��Ha�^s5+�s�ލ�j�U�\:�
� c=uI�R\ݏ��V�,�f���`� Iַ�_�ͷ�$m���r�F)��5H_05͵�ɳ���m1n5�!:7�OFګl.�rqW{,J?"g`�v�qF�z�B�hAb�~�%k����@�����p�9���F9��MhJ�JtN╨�v~�����Քs^!Z��a�ظc/��J��~�"�aeiևLP�;5Q�x򛒧Cǘ�ؓ�2q)Ţ�un������)H�9zJ1)f/qo�K���,��.����:M[Q�Ȅ�����uM�}2U�е������#Q��Ë�E�7w�	��߇���(�yܖ�;��6 �,�mD���|�X|�R�s9�G�&�w��O�a��P�����RS{=�$U,����9<dĜq(z����YD�9�V�̧���\U�F���<���`�j/��_u$�)˦���pT��7��Q� yt=��h6��ڀ3�F^���T+�!�gi/�	�X�-Mo&u�`��`ә�pŴj���F�u6=�B=$�v��#	��_6�{Ǒ�Z��AH�P��,�[����M�Ql�/�[' �-z�p����:�4��}FC�~������P�V7� ZT6}�<�s�D�[Ť,qX2U�$iʚ���81Z�N�hq)�ei�P	�C�;'�x���qG�jc�0#��|������=H-o���^9�\朌x/�U^����.��>c;_`8�Lwʂɉ7��#�~���U���f�o)��#�2)e���N*S�uE%{�F `��Ì��N�T�,C��{�N�X�f����7��n����;�����q=��mF�/����5;��ٕ��Ҟm����+l~��^��������o��5����8e���;L3�qA��� �Gp����e!�-�>1�؜kɔB8j�&b6ɑ���_����{(���c�֕��̨�]vh�e*�W/{��b4�ߑ�2�ё���=������3���R�k�☒�� +��A F,��7dl��%:S	I���X� ���G����^ �@�5���o���Rm}k�m��M�U��@�P�qyF����b$�Օ��D�x{��!���(�)`����="f\�7��E@�T<b+�)�<�t�z:�����ݞ��h�p��ͺ��I�v��}���v������F��s>睽Èl��h�X(���F�V�R��!�&m--+��#���rѨ^[��QjYO��>�gj�V���$��ج)N�t>��,�;P��^G�ޚ�&�{���ymy='v�/�&s[n�2�gρ$f��=�V�>���}����v��Mԇ����,�5a���I�C��FL�SY oh�"��e�6�t�s6�\�U�輇��U�����n���h6Yw�A�ƥ��͉%�N=J��%���B�6e�lx��L�k$խ��#�*e����}P!%8QLg��T	�D���v+���ǐy��]a��T�@*4�y0C���U~9\����b1�WQ���%�����=��و%2J��2����y�/Ce]������1-��� ��J{�Ɨ�cn)Č���榱r
u[1�_Iڶ���Q#�jjCrd7������.Ƞ�eo��D�,d*���&X�[4�HBΜ�&H�?����ph*��z!��Ԛ5Ff[Sm�9��/��PbL�m���	(y	�Vڰm�s_A�H`��3 �OP�F��gU%���e/����%��rP&��>�z �^��ck����Ǚ�����ְN��R�)�.��IP^v�L`#��1 ayq��V%���Q�u�҄@xU�M���pE`lũ�[R�
��2^8��2y��L2K�j�H�Ӻ|���x{[����7?]`Ҫ�9}����#�Pѫ��`����R����'�nK���TL$R������z���i�`���HJ:��q�+��F��z������z������6J\��.s J��H6�wZ�R��B]��0d.�WM)�=G�
xi�<?����(����~�HQ��䶫��6���������,%�4ݝ�3o�5��}
q����W��*rHZ�����T�O��������I�oz]J�十<�}w@q:��k�.:�B;���:/#H��N�/2i��	�L�6��������V~ï��YCݵ������]WQA`�,a��@P�]N79B���z�%�!J�O��m|o���S�U�Φ�4,Y�����a(䛸yx��M��銖ZD�|�m�C+�VqG#��x6]p��$T��)�ʙ� M��f>O��	TQ���������+�C��bX<�C�\^����{F���}���ޒ�`�Vah����p�˅�Æ�{^!�λg�(��}P]��� ��c,l'��s0��!�id.d'sq�F�oCL�-�k�9�+bX##��d�H�n�G���#M�ŋѴf�v]wv��F�]��jP\�<X�y=,\���'8F[�A�_A�mqE��Nl����4���7�Y��n]�b;��7��{j�fk<ܓ]k�F���`�_�V�����c�1��=/N][ΓΐK��Ds!o��k~N��@!�l' ��V�L�?�������[�R �raM��ϐ�T���������S!��h���;��Kֹ��-l�&�� GO����	�����,���Ƈ.�+L����7r�$c��ք����!��Y��yt� M��e *�ϛ�xs[Q�T�
���!3F{��喧NxR����.1��6pbcw�}xnT�y�{g����$;2S�U��Q�ÉU������A�5
9�q;ӗ�?���;=;���	���t����T��H'< 
���j�t�&����§���g�B�
`Y����G�W�>ӎ0W�;Q����!������N�'����dw�����.{��`%��2w�H��f�X�~fP��M(�	�lw���������R�D���M�8�����i�=�%��b1J�ʕ�/��.�����Ay��dE]Ks�'�D#������j�����
ױ�T�՘���|���0��v���$�����"��!lo�$N��S�: hI����սmw��/�5���9�]>�"�����xEx�Kp�ĨK�9�RT�.�����-���->ٝ��7!W�6 b��/�n$s���^c����y�r���'A@�x��.��D��{���`��h�G�t�j�e#b��t���া��,��(e^�v�8QI��]�=�e�[����h�_��8e�M���z����*&�Ozs�2-�!J.�L�b��-'�
A���U���U�e9B�ܔ{�y!6D����0�>�*�z�0��j�!!q^`}�'�=3f"��C �2�8��nr�����2`�r�*/����T���^��*ˇ��ĆQ:��Q�y���zC�zb�-�;_Ҋ�Q)^"?�m^v���)�,���{ѹ7p��򴲏�p��*7YJ�����E��g��<Ez��#]�B�:[t����&�Mc⚫iƼ��贩?EƑE�e=�'�+@�!�8��FG&�oś^7�@g��xΚ~�#����7��)օ١�B6\�ݓ8קߋy�/��ק�M^%����#����<�_�o����F�tMB_�@W���.W��D�
t�>8ᰫ��php���x5�����/5�?!k�i�doǁ�Ŵ�bE�S�&�c����J�>�<�����r�%��i��7��}�5��V����H�����T����)n���q�������:̮󊰤��d^r�~�暒D�<��*AXa�_����: �o���լ9eT�Z;��Fk_�N�=��sĜ���O�שƷU�����K���Њ8bh9�u�Њw�(�޷�*����q��ߊ4��Go��R��>S�[k����G�3$��5�u�� �`,�T�ӗ���}T�8un΄��¡$	�y�.���f'��.5K<�w������מ*���*��:V�j.酟3�)�y���Mh� ��*3�m�}n|��_�P��	b�?� ���������#�W8�@��|���@�*\.��]_�3T�W3�]�0L���i� ��bhY�`I���z@����w�SIy������x��k����ii����#�r�}�d9�%��El:�c�~���0O���� z�,/_.�|K"���$�(�_;)u�>|҅`m� �����U��h���v�!�<Jμ�"�Y5�� �X��,'p��8��B�v�C]f|��������9�cy�,��5��VC�z��N�5�m3� �W���Y���ի�Y5C�="L����*;�X�&�(K8��t�i�]�^�ҙo�KJ���)�1����|m'p�ع
X�û�nn���kS�oC��J�@����F�F����iM>��x�m�����Z��{*��j¥���^��^����D-?F��]:uH1}E$��&f���Ǵ��!��S]ы�<0���m�r'.@�� ���^�jvv<*LGɈ�L|�,�+z�3j:��e� �qk8�\��`h��u� �yr�mf�x���j�L{��onc�<W�;��i\K���2ehI���Q��zb��6k�\^'��yiQ�ػ��;�5��	�F�TB�$��U����0{r��dӈr�Kn���ab*��*|J24�/kP�}
b�^�|���,�F�/b��'�������蔞0�#66M3�L9��.�!X�cQ��(o24>�����i�.w�w'AŸ��Q�A�)"ǩ�u�P(K��f2��M�(���[I*����Ҕ����{kXm3Rʦ��_��f&�<}��w*#�_>�aI��TӤNVl<�&KGU6Fkp�r��&n|eƪ��@`�,�r1��i�0���G
s��eGʵ����4�{���	��Bt���Ic�9\v���w��'i4|^>Q�n��*_�;������ϼ�@�"b�#�=L�	�@��.���tr�Z�)2�w��N5��R�Kև BmFܒ�0��A�Bam&�,�����Z�1ϫ|&龨㯟N>C�SG/��.6�D�V:�6��@q6�4߮.��
4p��c�³>��ӵ՟��t[t���y<D�Z9YO4�)K��8��w�>�����9�>�H�� �"�P|t�^>D>q3ٞ�c�B�N�������l(\�	86�4���*�v���/i����*g=^�hINř^
r})TK�*lR&ױ�!�U����Z�tt�#�s@��u|�j��F���d�O�b�9�7��t�X�q������\��79o�b�s83%|>sý@�x�.`�a)���W���X1(�1=]~C�w�Ζ>v�Xs�wכGO�Ճ�K�h�� �=���i66����'F{��+�H[�{-����ޅO�0�ȗb5PAo+�V<nV��]'Ȉ�HV~�p��*����V: �z\Ɔ;0�˵j�2�UmHD��\������W�~���X�uvBĶPB�;�X)�F>�9��t#�HFR��'z���w�fH��Z�[uF�+���p�,;5B�w:���:X��K����s�x��zN�D�H������2`��v���yذ[����tE�Z��ś�Q�[���n|!ލu9j>�����n��V$�t�F$��*�
͌�pz��=�Sÿ� ��v~ti�t��,5g�c�.�f5ԑAN�����*��f��]������AH����O�;����M��Zj�T��@�l2=�d�1��j?mgt��'J��]D�.
��`�W�¾^���y���޽}�l����,Y���I������L%A��]/�&0ruF�Y� X��#G����j��Ag��H}vxd.|+����Ь����Z���� Ѥmr�6b	��U�*u�|�����(NR �W|	Ӱv�2��݁�#'g\==-�g��	C*T��}�+��h�m�ͼF�SZ��SK��#�@B���I�pf����s�N��e��ob�d�%+�m������̖�FCc���'E�����d��W�2�:U�^�-t��NV�X�/!E��M:���YM��a��f������{ބDX�@���2�3�C5�&�(�5:�D"WRB�@�k2i��m>>�k���9=S����ߦ3�r�W&��h��!����%�=��]�C�}����L�<����]��Hߦ�>��!QQH$��)��hhGڕn�h%�`�-Z�i��+ufǻ��8J	hM�Ɔs�}@E���"�N�;u�2��ɿ�_)�҅�g�d�ޱ��X1`�SL�b����t��l��_CnA��;�'|=���τ�|ry�{�����mh�<��6i�$�<H�4������yD�;�UNY��R��p�@?�^�&�l��x�+���v�������ռƱv\1n}"g�#S�1���������
�CmI����z�#�9�d���d2/S� ���os�#��n6]�����j�f���Ɵ!�y��U�("���n��h7zh��)75 �olgU���(��S�
18���o����>�@��X���r~�4Կ����
���$�����6�3���j8� Rt;ܨ�'�]�9���h(4w�lфG���][5��*zfi�y��!�L��� ��j�ڲ�'����A
m��~*ND!D����GJ���h�@�PG�R�H��$���k�4���U����qV�;؅s}�Y���+U�o�U��� ��'Wb!���v,\4��t���lFv���,B3����A�pG���^9z�Ɛ��w�P��_�-�j�Rq@�Y>��"�\����&�0;����Q����kK�$C�{ i�&3����!���39�V��`�|��:s���f��C�v�S�;7�+]��)�Lr0l�ֺ�4k��6%&��!0���=U�@��(s��[]�Q�&���^�1���o�C�Q�fl8x;��2�yo/�#�޲��jcd���0����]N��Y��1����h����C��6}��������@��,�+I�ݠ�-��J�f|� r��+��j��?]2P��gKφ�j"��zq��A�	��n;XiKZ8Gs��5!V��ff�ݏR��w�Kؽ��$�0x)U�P�V/���4�s1�T(DД�V�%�q��jS�n�R�a�:���SP����w����+ǃ���c5�(��;��.�ɇI(���L(�<�f�8<f0��lKZ]Ѿ�Z�Ft�HB�ʓ��NF�{}Q��	E&i_R�,�1��uҟndO����f�Jյ'��*�/���1�_MH�ӭ����5��[RЎ���V�7�%�%c	�/+��M���9�F�O�U1;E�T%C�*&S�A��$�@!G�iD�OP��LRKgB�^�D�v������u��zsF0�8�
�uL�:%��$[)%���1?Y�Q�t������u��Ϻ��*G,#���G���rx�7�k�����Ѡ7�Nl��Z��ơ/A7;S�eI�;`�����$ �+���U},e�v��f9�x����>7(�L��T�V�O.�����bnR��R�o� X#���h�pm�
�I��h���/vA��P	��/"�9���o=����F�e�ݰ"z�SJ. ����J�k��ݷ����Hm���^����Z����̘�Z���vt4����N'��3�J�$���w�U<� -h�?B�!͠��P%�X��de:1��ȜM�5/|��+Α&^w-d�p���c�3����Y�X2�9���]?���~Gt�Q�z`3�|��[��I�\6Xw1?g��w����6{��4:4+:���e�D�л�vB���s<�~����ɓ�# �>�
8(�����BO�Q_ TBd�f�T*��|��T�!``K#��$wq�1\��){��{Uhg���_�@n>��
A��Y�F�7�?LE�[$�vi$5hDS�i[EKG%���[饣!u���,��]#�pn0�p�C��<d�p�ܝ!�>��v�����{���8X�0\~*R^ه:�9���{��d��!��1f_�B�mO�,�E�U�	��ZH��K�+��N�����������N��0��MBLZ��̩+!��	]]z8@H��M��7M�m��?J��L{@9�bT�t�?�H(c�n9R� ��O�mXϕ�� ���6/���������:[Y������[s�^�TX�S���k�$�&BRG�A߶ntc��6@��Y�̔������[g�v�R�>����Dl��AQ�-��rOg�d��r=;
�$)����xD�lM�T������k1ԛ�����Y�Ǚ
N��72�j��mё�
�t��1d\ą@��8(4��R{�ծ�盡�<σ���k�b׊k�޴~��	@٘O�^�Q��+MK=a���P�CY$�p����uD�dO�e�˕$��@�a�c� �տP������2f@y��ݼI��sW\\yp���b��G�wP;��Y�O�;R�2q�,
(ݤ�(��ǹY�=�����I$�������Dں�xC�7ZP^����t^-Nǋ�pw)�؎�b�R�X��r��Ś���%
t����!�~3F�e(�N�;��Q��ʑZc>�Y\��xv��S���g��3�>cC��U˨�T�G˃V���6���(���iǋ>[�>%o䚹������\`��_��^|��.� �(��Yvi�@F%#����h <Ҥ �H�y'�Au���NH(��f��?�g��n��R��'�sI�X}$��5�^�V悊����Yz9��G�X�)�h[�Љ��c<ɂ�=q�Ln�g���`;�P��>>�J�ih`����ƭ1?̻���#�L໣ri\�/z���k�"�4����2X!�@~�i�⊪��'ً~�����;'�F���R͎���k=���Ef�u�骹���DYz�A&��!�����y������c�T��;w���$Bq��j$��^3v9�ҩ��H|	�lQ?�L�3��1"��Y׻��f�`g�?󥚪f�qA����4���N�2~�F���og�Y��f�PFi}�r���l"k#�%�[Y��v\[U�6�,潺��"��V<a��:C\�Xv#�+%�9M���kn���I�.������#������=?`E��Y�U�C���G��Cϱ�>d��cBK�#�Е�7��G��>׾�_����X�J#��	����B:�cU���k'�%����&�j$�0*���}]�șɭ�@Q}lxu)l4�N�$J-[8�)��M8R�^�cX{�է��ɛ
l���S!�9Ŋ�B"V����x�G�$�i��Gv����TZHO�ke;w��/�rU�%�{�*G51_���/H�Y��5��Kj�Rk��>���_a,߸@�_���/�O�ڃ�d3����j���_�(U�K���pR���p�\}݃#n v|`���U���>=��\��J�mDJ��V�3��YQ���������4ߪ&���@?0{�Db��,�l/hs�����B����S��J�F�L�A��}���ٳ�Gb�����{���m �%����5�ǩ��q�����L�#�"eK�Ό��t���RcSN�EƃA!/�>0�g��^ӌ��6-bUE#1�����"��@	;���7f)Cy��p~Z�#�$d��U>F�����z�t:�D����Yg�ٽ�F��,GKNf�_$T�y���(�>s�����i���6���ʞ��ǭ��R��&v�b����^ڠ�4��u�����#��������^O��n4�.�V��<ϲ��Ƹ�)��&��;U gܨ'�#%�Iر�M���%��V7IS�5˸�O�E����{�lg{�R-*��<�?���TX�#ߣ�e
pH,�t1��`(Yeަ�$�UP�)3ڿ^ {f�Ȑ�C�V����w�ۧK�Dl\V�G#9.rL�Nx@�I�ș���#���7�'����|�UϮ��0���-י\���9c�ȹ���.�#���Ye�[]6�'��)�(�gR�8 �5}��]XÊ"�� ��{*�W�j�(@401�bB"!6��ȍ���s��1����aT8�utHq*����Da�3�tw���e1�@e�Yo��ܘ�o4%�ҹ��H�+�Wչ�Fb�|S�Jk3������mx%�B�T��g�	lʽ��;�?�%?�k������n�*La��k,�@A�A���Yp�B��N�֞�����'���r9Ը�HW�y^��{)1X�ˡv��=Q��4^�:b�Y|~	�%Z	�[��TR.>�x,����%%X*ž�!��`��*Yg��_���E1�R�4��@�s����U��p̠'�� R-����n'$��V�´�Kwĥ���G.�[7�ҰJ���.��O
�(:8��Z1����� "�C	ȥ�e/�Fc�{�R$��H,�m���8D4��R��Fbq�~%4�%ݹ�4C�[��i�
�[��4Kx%� &�<�E��>������S��[s��$� ūF,,x;���%���B� �������<�����fƲ���Y:ד9y<I�����	M�NpI����#�$_X�R'y�fM&Z)�!QX���K4�o�̷U_n�b�v?yX� W|EW��7��H��;�E�H�n��)+��pͱ���GJ�?2�tg���y�XU�ѳa��ܧC�(nQm�[m�<��2��@�Nq(�Ϳ-����|��}���y�W��!��'�#�3�|�3�ɏ�%�쀟��o�w�R8�H�榛I����3{��NN����MTa��>)M�jvݯ�V��(�GF[������> T ����[3V�@���3<��TLw�O�Jq��Q�Q�p#�3�s���ʆD]��&٧`��{n��i$�s$����#��$�ռm}L�P�@T�'G�5V��[p�_������n�E�U� �С�f��I������ˉ���]r/@��TQ�=,��9 �WV�i�v�!��b�-����j����pg���"�X��p�vӸ�v�z,ɍbTʀŲM[z��G]�L"���-��+���^��
�ѫ�u��T��@�a%
3�w�AV�C��UjM�g�a�@�zA0��h����X��%�N�D�5�w�<�ƴGk#)$tD�0���Tj���Da/��h��׋����0���ה�d�V�j�*_��ok|�ۧ���vx��K�/!���� "�h��<�[j;޿�>��?f��?����e��y���P�������:le�Q^�fI�¤��i\�9�eD6^���z�j��(���F{#P�$�_ͤ���1�fC�z��u
��>K��Ԩ��-�)ӎ�����1�]û�+�J*�b�z㠸5�:�MoW��u�&ʊ�@��ޞu,�`X.��q�z�ptC�"!(.Qzܘ����ђ���C�D��ĵ Z��X�O8�-�ȼ�`&.���t�T�Ɯ�\yXH8oH��3�)1Zj�=�hks�Ck^��O���#�h���^��#*U5C)�h@�:Z�}������v��;������5�QRp#���ԗ)�����wm����bQ�d�<���6�2��Y窷�⦁��t�uK���)b�߹?]�-��1Իq� Øjg��\�xp��(Є*GD��D��u�e�2Fܖq<ȝ�r�Cj:Յ�V��[���H��A�c)٨4���۱`̢��0yaѩ�N�	nmI=PJ����%��q�t�t��V�y���랋Ѝ̏K�{�|M�QK�G0�����z�%і����R��)���&����1Q�W��/>I�ҝc�%��bG[}c �婌��Z)���Q5٠���������OV ��[�%��Ӫy�!�
��$��]��N�����n=n��Y��s2vy�f�V�D�$��K���F���ߗ�Ai�ʻ���Ȯ)�D��2I3s����'?�}�g2��� HLD����>-��5>7��c���7�-�n-=���%��9��'�j_�Q�?P����<����jLs�ڛN
�	w��ac����s�m����Ʉ���P�
�9' ��k��)��M���3�"r�8Ρ[�[����57�,��,�Q�=̞�n
�Ի�T�7a�?z��V��/2�5 �^�&ԇ�`��|t���l7B�kJ!��t�⃒"T
w���#Z*C�%��'�O4J����6�M,-@O9�*d�����bxg,�?��
��^������-̿'Y ��"�M�80�9�{������n�D��$�F�ϔr���@�����XsPO{�iT��ƺ^�
j��	�tу�ip5���}���q>na�o�@�Ic@����N3g��oJ�jx�4��.��a�D>%���~��?p�� ��:�kN�m�ȌAt߂8:��=8Kׁ�TbI�*,� ����|f�<��)���i�/����K��|�,�+ۆs��J��|�4�
Y�4&1��
B��#��<��p��A��觖u:X&l�j7*Q����8���2laם�.0��+���Q;s�\A&� ���◓�lЀ��?W�T��$d#!U��&�������Q՗Փ�B;r��jX�SYd���~��x��:ƈQ�缩>5�����nl5�^��J�kz�1 G�X����Dx�}`V��p���WS�HP�n,Pw���i»�HDS�hG�xכV���I��)p�K��˻G3΅"Bq�PS�u�L��`�$�nYu�LZ'���u��\@���#gOL�Z@(���, A��㦬rEu�[���}X�,Sn&�&ĺ!��Ϊq�ƶ�ٲ�Q_�����G�j�k��Ո;�@˹�|G�yd�`����?:�>}�g5�M�5%i,��]�P�0֑+�:�(��Տ���N��&^�ɶH��ne<VN@b�lw�=����Q[���%�G�V8���j��M�:Rk�AŤ`P&�SD�9,�S�[_ }N��Ve&����uS,��Z�s5��J��`9W��7��ҏ��jF��-����4�l�)�k
��7\;��T��-�p���@�'e��i)�]_���� �ge0 ~�{V��n�J���Џ���d1�����S6��hg�k08c#�ǃ��ZYZ�1�v�l��ÐyYZ�;�'9�WK@NN����;��U�>BF�پ�!�t0�6�LZ�o�T���i�`�E��e��SS���?oes�z��4���Ϥ �� �ν?,����}������WE~!T[r+�� ^V�ì�6�1+{%�~�S��j�
�`�3utMKs���*C��+�G�e1����1��&��Cs��!�|����Jq]i�<<���!>]�d9J��I�8)M;��Og�����,�+���P����[��G�}��^���$�[f�ݍ[�O�	F�R��*�Ӧ��1'��)����7G�nX�/�F�O���;�?���``"������a��Q<����7����JarV)U���p�R�z�	����,��B�@,�"iX%C�/Ѽ|y�Ȅ�9\�,����z�S�LP��E๨��R+u#	U�cE���JOy*3���΍V-��N�����M�I�s�@��
7N�z��x�}WU�Z�+�iM�z#t��OQ�Glj���)� ��qV�#��aωk���Ȓ	}rC"�
���8+��hя�W�!�6��F/9K���-g���#cy���ˑ<
e/SDK��Y=�&���:����.գM�mB���d���������$4��ws�EP��q��c&.�&6���>�7qx��H�tM	�!�|;?��@R����T��~c������6�0tw"(�V�l���}�0ѫ�܂���L�Z�V-	�)�&�M):���t�*��$�Oa�~�wu�� /LD��Is�k@��jȦY�ύ��>���L��'�5T�d/ء����(���[Ք�;Ic�S��2ǽ�gy(/��3Q�|j��7E���a|����&�����Ӳ�|O ��7q�N��#�u����}����#t�O��<�o�bt�	g}?V����*�q`�����l��|2Km��rx�H훯�>�Vh�W�*H�����G��vY������ۆ��YJ�#:H�[-�k�a�K�^��Vk�5p';������)L�&�^��G�6{�����gʄi�6�N�zq�6��ܟ����փ�۔h�� \�P�$�QU��{SzcF�h,�]c�f8�}dDζz�(��n�"�_Y��h�+n�[��r�����
aw�v�T2����g��H�����׬��������<�_���]�����.d��C��J�����8�qT�ɠ�uֱ���0F�����rB�g8�&vd�B�Q�s?������1�}KԩRCv�&��/	[���Pp������'M�zb���ʬz �I2�����V2�����f�;\G���9�M��t���MD?W�_e�g��pv�kȪ���w�
�t?6v�ht�� A`S��tO�+�F��*�!��5��ٱ�*��y�!_ߜځDpM���
����X���e�C?�E"��@��>�4*�"������'���&��[�O�����wϻj�2>������q��>f單Q �<ls�_��KSGV7V�G{B��̝�qoJ�si+��'�!ջD������Q�[X���j%�J��[�-��"�J�n�R�8��*�b~P>�����{27e���W���?��N��~���)��y
�&����� ^5���U��O+x��gp���oT-�[q=E\�7��}/�q�o��-��Y�� ]�P*)����,�D��w�Ә9quM�!�5]:Ǻ��VZ������|i���˫1�$�7������bs}8.^���׫7h`���"
mCX�+ s|L��~;��C<(��Yu�_��J�HІ���?�;���_f�*���@n>�0�Me�w��X��w����]\k�K7n��ڊD�����(:���ؚ�o�n��u30�[`��\Gx�����=):�D^m��	W�է��o�rgĒܹoyhYƲ�<�%1����F�����s��DVss����bV_-4?I�v�hb�Y{ϑq�v|%�N;�s�3�nn������BD٩ �^������Ԧ��H��c�-�і�)���M5��_}��ٱ>L04��� K >��C�� z�u)x1����i��f�����V3�e�k|mip��q��j��e��қ�#Z]�*�zc��
�D�KP?��OI�*r�vK'����n��㬬���X�\v�~;��3�o/·<�I���Og_��rv�c}�v�H�9�OcPn���XԨW��a=���`�3�p#�+� `��-�_6G��	�R�K?B����x�!q��G�
^=2X��0�Kߕ;�����<8C�I6��l���d.��!H�H�D�>���G2�6���U��l�lv�?=����fq�9�[�F�n���6'|�;�3��-2��X�4��eʂV��@P�	�\���^]�e2����!�9)i���, ��*&j�F[�ӟ�!iVR��ɯ��p$�����x�y
�)����֥.���8#��y���~��\��mR�t��t��ծ�F:~�4���K�R�;<b�edB �֚Or�\Ӟ犩���EuV�Z��+DC���}�9��bɄ�^�R�W}\.�T˖7��q�=�҇�����4��FmUJ�t� �!��*�_L��rJ�Ą�D)���ؙ�$PGB�/�6��7|�p������4&0K��:'�rx@xc����(e,��>��od�2[�b@j�j�xo1H�{�������Md�@��X��tv�PƜz|��U&�Z:��fLd�1��Y�Q燺 �R�-Us1����7�q&h�MZ�@k&��	U��+�8A�T�ue�ȡ���'�:{UY�H�=�b��p��nh����M��rv�w���Dܷ�����}"C��_�?��0���.D�)*D[Ԁ���@�������\���h؏mȗd�G�&�����H�IW�ɕM�$�D� I
u��^u����&�o3�݊|�wӃb��/�A<nC�޽��&	�yx	��W
��}mυ6uf[�&��U$���H��^�� �p����=�;�O���X�h�	4}`�X�6�]���}��֜���U�H	��Z,��Cr����Cc.�kF��(3޵K�b���m��*���D�p�c��\Ukć,XC��|P�Hā�݂���GY��N��x>�D���z�u�r�<J�O�� �ź���ݒU����p����C��:�7���A=�J�/(�����q�w���%lMYq��B��5�I�9-�9�!Q�u��5I��r�����6���芇ԑ`pi��H���t��tߎ<F��m"���u6�T,ج�kăc7����&���/sA���I&||�P�����'�rj�eoaZY�Va�W�:%�f�H��I��t�KM&�c��� �,Õ��_��X]vv�.��h��WCe��]{^?Ûh��U��a_	�ɞ:O��8�C��r/a#�xD��n�����iJ�x��Li������1N�{DO�/-:�{�5�I�������qi�����U1�~�N>T���l�ّp1IC5�8O�o�T�@(L����=.m�5���1�.��<j9�T>I/�;+��|�b���
1{^?ȣ���k�%�ݵ�2�ܨ�r��;+���T试�5v����
��G輲�a.@��E��G)��2<�qJ�$� �T�Z!�X�:P���p_��!C�䙴�CAw��@=
���`<"���	�a��b=�d jiT���>f�?1�?\�s�o.y�񒏣��AG�>*�G��nP(I}|Xwx,�F�����X2ݥ3H��JF
S�gH.i!�6����W���s�y�|��PQ�>:�H�c�)/�����"$![�F���|]���g.��(�,��T�~�-�!%#@@��6'�͟������-N]������,�W{��6��P��M@�qk�=��-��Vkf0�e[��5��3�2j�4{�������s�y¦̆�$ٍ���.���[�h�S�G䰙Y���~� K���2��1�&GLv�xw=��oBT�{�^3 /&#��!nB�et�E	��<���}z	YlM�Ɓհ���W�/��];\�M$Ý��|���R�T�lb�$XЇLDc?��V�