��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&��n?��1ů��> K�-� �&�T�Ek/ֆ�\�놭5�DꢘP���+L+X�4��J��#�0�8���������l��jT��+�(���������6�MC!D�;�m�퓊D@v_p��䙋ⲝ��C_�6�Ռ��#�� ���	RD�4D��畓7���vn�H���0���fX����4 �CS�C`{��;�L����li��� y+����FD�p"��]���y��R��K�({� .؜M�������	^5���ɋ��&���&�@*���
e�� �t+���
_6��O<��7f�M��u���m(MrN����z�jL���@T`��M3��c�uQ�Y���%�dD���,�~^���y@Ga��(����C����	��G�86�S$��ɳT�ز8���:r��/y�[ݦڍ#A�����i�&<nU��<[5)�Z�-Ĭv���0t���d���"_���:�'-��d��*��q����_d�y�N-��~";#��������Y��؆���	6ZJnԷW��έ$Y�K�?�4���L�w�Wmiɶ��Y�?jx#*�i���F�m�E����O6T>]i�_�9;�!(��kH7�OS��_��[-M�((��lO�s�$�g�x7`��ZV�E���F��,9�j	@���]}<�ahb5~ãdl&I^�	v����-�@�@���	��!��d��`j[Q��� r��;f�i�.�m+UH7��/OV��c��������l��i��M��*'��?���G� SK�M��H?�ç��q;��)��Rȩ�"@���r��Ml>8!�S��L��EgeH]�8��>]GR=&���C��i�Za�z�,�F��h�q��^���wT�a���%�9�n��?~SИſ~�mu�OlIv�4'sT���/a��^��9��*��G�Fh�DM�_��CN�<�_Pg��O5��}s�%��m�o߫R���X�Q?��dK�Z|:�=��y�P�)���o/�d\�6�� .���GJ���tՕ3)��D�6�Oj � ���b|�Q�ϜkY+\1aM�h�T�y�Ӂ:���$�2��D1C����]�SY�H���Y3c�CJ��H�>����jꏵ�[3��ˈ|��$
GU	�m!W�������+t&�9�O!�%뤓*m��:?	Kgix��ف���x��x>�ދE�M�r�%�\n�a/��m�`y1w���{-:S*@K��AW�T)�jԹ ҃�RkV����b!�⾠u㾒���$���<z����>;���i���6.���6���b�!r���P�y
�.a6�+L�
_t:"��ɤ�إ�&y�*��ey��;�і���Z�y&�a�uC��,B�Cn����eO~����d�I�s�����ɭ=
��M;d@���6x�7��+]����Zc�k|#�eVv�Q΍Emtm4�@[�����k�\���Y꺡㝗o��g��?<i:�Sw�N�[4�)���LdV�����9���C�|���#�Zj`� �`v�T��ۙj�@1��R��pq����L����z1~���Յ���~K�ă�6���m��qGC�'�� �L�����4����uw$r�d
{�V�'�[G�9 �(]��n;4���-���Y�����La,.���<I��]iAI��v����JҦ�u��Ey�͈cWF��� <*BZ��Z4�������J�+J��i�JI �s�rB�,Q�7P_qrq�@L�fXM���w��j˙���v��CS�H��I1�?� �)��0}�;Ք�3a�d��ܼE0ROfJK�b�6��������K3��i|�JG3���T��qʽ'N{�δX�Ao���:��X�WטS�|�۵-Lh)�/�(�3>��6��ܳ�|4��$H�ȍ^E0
�4�A��G��r��w�Pk7�W�Զ']�ֶ�:�u
k�q�� ���`e�ʳ�\11-�8$�x��uS�k0�/�wo�!t�\���)w�k��$����8��EWv��������
�EL���pZ�W'�&`A(LO83�E�҉s;W�	z�٫YJ�y3k��+��N9(�D�t�H��W��f1C���3�2�u���w��{��v)�}�܌�R���`ŗ��W�Yh�ìkhc�v'FED�x�\�a8���8$wǉa��+���B��HZ�Lii�/
95@w�޲�ݧf���[�������줊�|m�#B�b[�q���e���M{{P9�t��0L�,l�ڭ�x$<]��bf�k�;K#_��`���2�H������9��"s��y*e�ҩo��ȁ�	3���G�;Ë���;7x&;���aS�H���!}.T%��əvL:-y�1����*���� �(�KQ���Qc2����I������Е(��3*)��x�����8M=�"Z��D���D�T��]̑#p�~�C��+���o��I��H�j�i%a}��5�����S*�����#J�.d'7&:�<��L���v��Fwn!�E�2y��֬ˠUj���J�&��?:qǩ�����|�E<�(�T�anE$��31�����}+?}]�G����7ys�*�$��q���iZ���gh�t�y���0:8���fk�ɤZB��H�A�_�<#/�y�E�J
v"&�qW�S�q"?�{MI�Z�[��S��P-y��P�?~�I�2��U�~��qfb�[t��B ?�{�h����ܵ���r�p~�+���"üW��u�W�˦�sW&�#W?�9Y��J^6Y?'`őFYlD��9�g9��S<�c��)bi/���#�+�/�w6'y1���+cê����qb,-}E&S��,D�A��ӏ���@���Pz�[_ύ��M��.�>Ѓ���sS5��)G��\ҥ�!�l�-�����b��e�����}��r�,�GY���U��`�[Ѭ̛k�j�X� �zIp_�	�)n��&�:�߭�.B1�	�G͖f��;� F-S��@���Ir	;H���}�Is0�^}��V�d���E��"�𶹇u��_(	5*�IN�w�3������� 2�;�f�ʮ��W�s2���D⑨`w�9�F~8;�!����=�p�6z|����o>�"야��J�*j$�������Is!�ʅ5��Qt3��۹��|�9 f��t`������v� u�ѣ(����%뢴-j
Q�;}��7�$�˙ּ�B��	��9A"Fr�\qrȓ��>�=�t�K�	���4��1蹖8��r"�\��&k�s���M���s~5)�+D��Rl%�`*0{@I�''���wž��}8��}N�0�@^�1��[:�� �|��mrp!d��TZ������{h�ɣ'�������yC�8��$nA� .Z%-�_q��u+����{~H��o$^��!�쀆u�W2� �
JD������)�*lծZp�F��x�%��"��d�W�V�_��x��P�/���a�H丐g���OVi�F
qI�]����'�9f7����B�i;챼2e���AL����&_�����Uǟ60��m}����+l9�+��9_\v�Q���Ust������_����<����GB��)�S]�ߤͺ�är�J�ѥ�pf��o,�5��U���߈ @ ��V�,��,ۉ�h�An�|;r�P��*1�b�2�+��uO 	�[=z���3�T���9m�m�
���ׄn1hx���95{o���9�w������7�SVՍ�awB�����m�3#�2�J1��������}��9�X�� �{��9JEq�㢉a��H�1�G�B�\��j�R�t�=�;.ޏr�޸b۪�W[Qz���s�+�&H���9�W��!u�cv�D�ɸ* �#�x-n/sv� ��g�w�Zp��7_k�����d,�$����mu�v�)�9mHm�	�Pw%�g~�8o�ϰ ��XL'*�BnMd��no�% o+7.�,؛"�ffߢ�s
�\.��L��M�n�E��1����ޘ�Pg9�X���+��ú�⠯�UZ�8i[����|+�:���wVV�.F/3��)]�SJ�PJz"�@��������ȭX�v!P$�P��MW��R���s<��U��D�a^�i*�*��*��z�fo9�mLE���E`�V�˦��0B���d�� ��7$����x>�r����8��W�����w���P�n 7d�f�ǥ��B����-5=�39��n�)�T��������1�3i}:�-#?��6�!�D٨�)�H2x����hА��F�L�b�l#`���q6:����R���t��,�B+h%�{c��
��Wg��I�柸��^��*��|�e]n8�=#��n2�2�|*�Fh�ۇ�T�	�l��d$A������?����=��ۻ�o������"x����`�0�qb\F긝RrV\+J�m��bfj;�
�Q e�7�6��T�Dj�7f�<��:[�:-D�ʄ�e�Jz�O�/����8���mXSo;��[c\	NX{���
{oe::*D�֡4���/ �~�7]}�	(˳�����cd�m��"��W��'��y)�>_F��P:G/VE�3a�h�~�G� ��x~g7���#�$;�x�L�[�ܪ`�D�eq��Ǜ����Z��.����&sY�$��Od@8�V�P��]���0�[:d�����wS�ӄ�6�n떚�,L~��'i�2	Z�Q&�0%[&V���[g�/�ǉ)�JXx�������'�5�����\ԨDl$Q��e�6��ϣ�n<���~lqHt<�����簴�o�Do�G݂o8ǿާ�$4�{�W���VC����^*u�kG��XJ����ʸ(�I�]�'p���..���M�ub�̡(U��@5�d%�����)�^����27��@��h�&H�+QtW��Hy�V�6r�lÕ��L@��P�9xP��Ɋ����{���Ϛ%9��O+��G�#����MIzh��7~.�@�L�)O��`���z�/������2�*]��08Wj�D�X���i]�o�+�%5�G�V�qm�'�n��� �B�g���x~�R�v�g�0ǹ�vU�".��	iD��֫��i�x5+C��?�.�k��ǥo|�:�!����f,�t�ㄲ��y�Ɣ�0��edU�.�y��C��-���^oW����q�Yg��/��@�?	n�	�D�z|�\%�iF�,u�0�Mm�^Z�ҝ�8g���Q�^jW�AMc���55�v%AmU�UHX	��R��@t����|�>Ԗ�	���w�N�!3�A��I�j&M9�}�h"c����Dm�i
�Q\֯����~�+��*+f��6��\�Q��㦋-�N�?ſ(qoV��[V�Ʊ����0�(Y�[��%[��iq��2��c���C�/Ԥ��i�QYX�t&��5B��\�Dm�ڨ9��?	s����љ'h�C7#o4�AY��CTe�C��5}�PoȊ�������Y	ڹ��(�y����mY�Y��%K�^����a��B�����K�X*c�'��.ᛙ��{���q��Y���_&�H�b��S%�;��(�g%۹vЋ���bo( �{`����*V�܋I���S ������M�^�1&`ˤm��i,˾�ls�� Q�)�h�|��knͰ�P���n<�,}T>�?��O_��(s<�����>.K��ݪ��j�y�����ׯ�~�A�D��a�N�I?Ar�=��x-@�zx��.�U��A�ZR�[����^��h.l�fU ����M�:N��O��a��8�n�5��C�t��Q��,P����׀�UR��+'i^�Kd��^_�X�Q>^��f3O�܂�*`�����R��˜g8����	nP�a⦌_l|�XD޸�`���a$j�6��_"M��n��{��a��6��zGhå��#�5�)��aʩ^�S�@�t�p��);�\�!�D��NH8�����?���ND�k�[�~��n�"�b�¢���Mqŷ	Jzm��͕	��;��z>�q��v��(�v�ce�2E� f�Ś�����h_�����F�x�d�>1���ZE^װ�}�TǋN���ǜ��6�.Ӎ������L����x��p-:��[�F�]%��tM=)`s(Z���0�P܉�;�`&̽_�t���m<�&��*�����ڹϯ��jꭱU�)�B��m#���L�*c|?YZUj����ϧ��G����AÀ�sa\I�\Ef�jZ�~�f�1�?1�W��=: �`d�C{ :��^$c	^K��xD�N\��Cgw�d��>G����:��Gxy�����k�"ӆj³���J\* J��)#.���3V���n�L����(}�F��<&�P�o���u�ESR%���z�()j��05C�c���*�#����_;�偪i��)U+f&3����TW��{$Su ��R,[DJ.�Ii�4(1� B���׌�>L��x�[���uIŋ,x�;��F��E!u3�c  $�
��@G�<\"����-�l����w��?�� ӥR��t?&��d%k��Y�6�q�R����V_�'�&�n	��1bR�<ZM|8ykU�?(�MY6�N��Q_'�y��.%
�����IL��c��FB�`�]3~���B�9T���Zg� �K4k��M��R:�ƾ��ѽ�<.���ҕ��z_�c� J��}p�ei��^�%�Baj�5�����$�ws7@��涝��?����e�Cg�C ���_���&����T3(jgzO�>�ǣŤ���t�y!��:.���;K%3;�]�"h���:̚{r<ʢ[�ʉʩ�o�g��xF�����U����Kz�bGq]��M&��.�g���,j���fG�!,"��.���22��/�ީ)�Tt��S���63���v��=!\2��J5����oi�(!�Lx�^]WQ�����v���~	�἞��>�B�q����/�ǐ���~H�ҫ79 WC�W��}rW����h]�G*���Ma�Y��(��>[�����*r-�����X{3�j�i'����E��-�x<k���-���Q�hf{3΄��cU4��)\SZ�N�c)1��p&���\��Y"@�?��(��L��0Y:��ꤖ�3��ez���p7 ���o;Vg�bH�c�E�y�Z��%.�|��.@M�P��m����Z�5ri8LKR���QX�LBU<����O�=<Ji�+�^����21d�_q�E�P�������Hӭ�2��0���a]�ӖG�h��)V�>�|	©tҰ��,i����'e�lG�aQ�����q%��1�Hyã-i�<b�AiB sT昽�95��_��M�T��JzJu:h�3��r $����X����0x�8�yn���G�H�a݌�Q��-�����3��'���LA��j�L 7}[��|�~�F�{B�Ti���D��9ߖ��z�;����f@�PQ����@�0�%g���T+��9Q6?�U�JWV���Ӯ�'1$�vrxȴ�.���v}�f$��ܝ�At�x���`4 w /?�b{��H���������w��,�RS�J6��9�WZ��`l�_���mK!;82���?Xx��r��L�Hv���O�Z�)ԓ�mO������TQu��p�1���8�#	�*~�QS�і��_�*{|i���]���c�8�aQ�ۯ�+�����(@?� |e�ƞ ���-'d��~-�*�@"s8XP`].T�|@�ώ4�B�[=�=�y���G����pFZ��5�5;Q�*B��f�-&"����4O��xʼ.�{r4��Q�?eTGC����'!�oSw��|'#!S�u<j��O�^�l��j��q���Z&�<�o�2�ȯbSɶL3�;&8��G�2ʸ}M��
nq.�|�����u�'Sz�%�&#x�����Ud�g�[���z�C(7����[N�/�DbI݄﷑�;����gȔ�0_1�)�z�᠓^�2'� ;-5�ݫ��j���$_�_	_e�����f�$�?�`����u���^W��x��(k�Fh���<��Zb!x����(��R��C3�i"����5�C/:�v�$�?ҝ�RR�4J���:v�g7�����Q��JK�
��]�|�2�//�5�ikD���jO�>!��,v��(��������=cH�_�nq)��N
�F-6�k�)�[M;w)h�=ͮ5�S�G�3AN�s��r�.J�QHtT�$��+;���m��t��|�0��9��� ��(� �~��&�@#�WTRYT�MH~CC�<%��p��+|?�t���a�^�M��j�03��!ص��2�]��8'&ac\��Q��P/��������HڂwNC�d��\��5I����B��^�~�X~_�P�� Vv��}�ac�ɑ�9&��K;���'#%�y5�������V�F�?g�ܖݧ�Y|��{���r�o������f��h�D�;����O&��@Cd�����0��j�u����}%��P3���������G��-]�q�u�z؅��6ZL��UT+�6+t�ު�r�}q�������R_t�Vqz��c2��cJd��c��A$F�i�A�k�a��}*F>N,���lJ��F�6����qJU�ˎ1��$P���b:�=g�����M���s������$�n�2�a��2G%�q�Q�����S��[e�fe�ȱE�& }�?uU���I$-?����/�3%�,�kE����$��	@,\?��@�-p�ė:>������]w�)Z	�6���,�Ո�zt0;���`�E�� UD�ﬗ}O�H�}.�k�]�-�q#��P�lʳ6b.�z�í�����p�V~C�'J��?���jP���?&+=yx(���Ȼ;ey��g�̰��'�)1xM~
�5gx����¯fFNyW��Pn��bA��G����B�f�Ѝ#�Q>l�y�Җ�)|�?�)5�sS��Hcc�(C���rb���m�����w:����74�`$�W��<��(ׂ5���d^��m�|�Vr��i{+�hZB���<���+�U����4E0U��`䃂E�8s�j���}��p�&d�	v��l)�'J���(,�z��W��D��l~�\�*�IiL��*���"�;]���/�N�E2�N��s1_Z�(rh
O�6��e�\v��G0!�N�|�>��qoO�T|�χ)�,$>P=�,3h��b�+�ܧ�����5��"�un��K���2q��X�a�i�%\�{}V!�Y3?x�����Y��Ht������7��Y<��20w$9��d1E>�0�b�*�*��L0
4{��_2tu�Sn�Kiٺ�7g(>�&mե�Z��<�_r���l�M���Ȳ���ӓ.#�c1 P$��e1�����c^F���l���f�F�o��!�|u}:p��b�0�+<@S�G�D���s�>T���v��fN]Ol[��
�9bs�*{-��?��i,��&k��\��14CV�����y&1�k�1��^��sa����ݎ�Q;ă�uS-ɴ6����-uB���4��֠^�6��Ǵ:Ra�F�n��o&`�s���i�atf�p�@))*�9qT.m���u����8��-UɅ�4R���!d z@�,_�6-���\p�
垻�����:�@Sz2�7�},��{�����ĝ�v�ȶ���*��]�[�/��:(�zOfc�f�d@i�_B��솞�>���|D�w	��|��,�jփ'#Lb^���O�Mz^��>ꋗjy��y$����:�{x�wJ�>w�fs�1I�/J��p�	aZUk9 �����{�p����^��}@!Fէ9RtV(%Vm6��}C���7h7ye�ی\4�&���!s�G,!\9#5¸�e�W�S4H���3���V�� Zo��a�ө�!�0U7�E��p2��I� �u��dVĲ�蓟����$�R&s���-BVy�Z�?gu�CĠ?�ɬ�7h_�Nv�ǀ3��t}����K��K$�-�wB�zG��M��(T�<��mꗆPcu�Z��*GGW:��8pq?/��A�+2��((����������ZQe��m;
��~���\��(��|�@��@���۹u��Z ����XJqA/Z����_,��MY���;ӝy���#[·�ރ��
�>.�`���jl]����d�X���_C���.��B���� �B�F��������
����bO)ƴ^Ƶț�Z�d��,�-
kZ����?w��[�%S�V=�KF��ь�����VZu�Bњ".Э�>�@��|��o��J��PC��fcF*$�ݠj�y�P��&����^`�=e���DbF��5����5l���E��Ԇ>���B������%��6$\��}�\y�FB	.M��0�41n��_Is�K:i�,D�_ڼ��~���|%T���jy��
;Y��k!�f��5�p��z�{���;�+�g1I��]^rp��ԤI��tQ��q��k�m�k�/[c���ڴ�∄�}���h�nd��@$�l��kԪ�kSe�����c�w;�z��s�^N�L���-���#�,n�	��������9��ri�0��6�������*FZ������\���"Ȋ������ҁ��ВR�A�y�Z9�4�\"Yz2h���?�Ce�j��Up�CNY7�	�"���:��P�r����P�yQ�',��1E��?�t�$�) ��=�= S	��+_������c0�	*L�=�e�R���){�36��W��9����SZ����.�BiB?H��&R����d���R$(��xB\p%�����#x��_����5]^��:�h��\���Cí��|���͵X�K��$�����v���sȏ�3�. �_�q�6W�+��B�,%{�����6�����ij�}����.�z9�H��/eQ�4���,8*��E�2E��[��W�|�S���h���\�	=h*S�����	W���{4�ce?��|����.���g��2�c@�5�7 �8XtC��+���+m�ƟSs��f�S�k�
mg��t�0���w���ן�I��
$w�D
�^����[ɟ���}X����&F�9�)KL�G�E�2�n�WQ����5i�XŶ�tP9x���;A��"Ê��Ѻ~A�Abٛ�#:�~N��2��0j9����
������+�%���TN��_X�I�����z���.�| 嵋��a�&\�����ŲG��]�}EB�f��f0e�"]%���!���n�iQ�3���F���f0���5۹�ũ�hs�x�ZU~Q�� 
�h��)�{L3�qgL�W����1�3�"22�gh��g��H��|�rX޹�v�G�\�*]h`��THJ��ᮖf�?��_��N�Z�� _܇gz�QX0}�"�2��D���*��%g�={���x�MQ3�(��pR��rǺ�@xУ�ȽXi9�{Sn��(��$�;=y�Av
�W��w�	���1΃�@C�Y��;�w՗g���ޏ	�ڥ���[��9b6A�` �T�������|�-�y��(ώ���U;�\ z�y^����:`��(E�~�rs@�b/�,Qh�E7�|�yXE=si�Q2��w�F�p�	�~yҏ�W�����������m1<s>�%���x�<�B6���k{9>���2Ȕ�2�1Ó=�]��A�i�>��s�k^���Z�.�c��2���q��;�A>1Y7�
 ��~l�ag0���]|������0���a��UM2yƮrO\軭��"��ȷ[��E�������؎����#���=��H�j	'*�|�_��*���i�	w>�[>a��4���~�<�$e�QKYyé���jB�3�����4a`��Vx/u�kw��5�2y��%Y{��D
B�4	-ᢼ#�-t`�W��h8(	�mÑ�Q�j��'\�I�`[j3������T�t�
��EƅX��T-��L#� �_?䕒'�`ay�տ�{��ݢ�0b�k��B���� 9ސ/P��� ��k`�j��ڪ�����D�!�w���gh�+J�1x&��5�#��|�:���������PN��.����5SDFlv�9�Ϲ6'et! ]��6���V���.�
�2鼲(x45�P{�}�?HSq�$i�O�ޖ���z�!m��4� ��v0z�|�`�G��3��:~5ȉj�a���=��s�����4��2�/W9Fߣ�%�N܁��-��Y�lT�3��&ʠ�)�$V/%<����J�e��.?G�) eg%�a�*K���"f�}r�6!����s�,J�]7�<�z��l���zq�
I�*�Ŋ����=�8>@3���˻(���?��l�쀃�S)��v�Z	{8�O6s�7W��Sl5�VH���U7@i!F��f��h���e�r�Q��
s����[S6Kr
tuz����kY�j�M諨s�S�W��c������ig�@Ui���N?v�=e?v�7��uVȁ�
��b�^dv]����Cm2*m�H8$��u����*��LC��]�T�
��R�O�Գ�ʚ&�j�����0gԦ���`E�N:�2kf��>3LؑMm��j�	7���!�H��ev��km~B ���սH�l5�n�b�Kl6 �G�}a���37�1$85���-�fL��++M۬E�TD��o�F��h�^pu� �����7����n����)�g�����=L�0�˱nn�����VIqmg��j	'�����{��r�Q��"F&�1��-�2Xf4�$�&�y_
2 ���C��N1&E����P!�$�e�`=���k�`~��e߼���
o����d=ٶ��%���K?K��kEB���$���>_�"+�P�7(l��J�5H�J�����f
�ӯ/�� a�^�1X�3v��`h����O׀z��c�#}���ؒa�O���A=,�w���z:�Ag?k!��v�mn�f(0�'�9���M�^_B�#zW,���ȏ
e܍վJJ��V���D3����}tq�7��
K���+������в�u2��O+�e�L6L��y
wG�Q
/R��]&^���fXwO��.g�Â��o$ح�#%���+��8�m�)�a���%��E��7
ԈLT>�5�)�H��P2��]�o�����"={�I���`�Y�H��kgs#��嚁���]��,&�����߷�{Ѐ.�IĿ�%T���ࡇ���r�QU&�7.~�K;�W�5%��U�yL+eW��ݲ�(K�/Nh*,2�_�	>��\�
7R��߼a��E�L+��̥����M>i=Dǅ�hr�`����y�'lֲ���R?���K��}��Os�4g0ߢ�ڠ,����"�� �%zF�Q��=0��ngZ�}Q�����ȳ��'���=�:��.ѡQ�����eF���s�R���Kd�Gg TUF��E*G6�˵T#(�֎��;���nь�;�J��4�l�@)`I]>��J�s�����T����a�f7�K��]H�����ԏ���M&aF��Q���'�U�^L�[{84��8W"e�vv��F`g��ᡓ�@�� M˳�m�,XS��2�����_��\�#�X�\�l�@�"9�ݘ�|<%^��d,�L�i\9��$*{����	]Ȏn�K���]al�=�� ��k�;t��ٻ���Z����6�ox'��D�D�bR�>���W~ަ������}.�PJ���G��p��Lh�D�D��^��	(̗]��������s.M��sE 7�7�b��B���W��|��|�X�ﾑA}������[C2
��<��b��7R/b���;����M��#�}��KE1�D%��C����:��Q���0I'q;sb2�c�F�Q��q�δ���u8�dE���k�߻� �}�>�N�?i
w6���=������8+?��zbΆIo��˨�5=K�ZArN`���b<�"i{��OO( �M���t�U��]i���đ�U$S���D��)+�⬗n�7;�9 J#%B�N͆�!��mF\�^��ٴ��|wj�_�(���&E
�|KmlA��I˅Yb�Uҵ+#�b�I����N�c�o�D��~��s�8�;��<�F�����u���`䜈��S����"aC�NB��搯^�f+�{��+{o�{�����z�����rpw�2�L/C�R&�t�@�#Z��y.�__���M���KG�#�а�����z�ߌ�Z8�Z�7%���{��=�[������^9-��镊!|ۍ�X���U�@�E��_�J�ŊGf��I5�/�
�f�P �猵W������vO9N�|1���L�(^���J!����0��@�)7�>�1���Q{F��3{����s$��C����]4�I����7��*�n�n���)'�\��	��T��eQ�ԫ��̷�	5�e��Dc��֫�Iws������wgD��-��i���A����z(>�8�g*d3n*R.�(�I�{��-���tҊ"��O���|a�U�yD����~��%xTj�ۂP^��wqc��5�`

�� �ɲݥ��@��/,��n��VD^��;�����8��|����Bh���.��Pi��y�uY&xs�u��Sb-�������2؋	)l!/��8�'�FPw��̄ڑ�~�1�5n�,��Sj~�5��]�%x.6ƴ���k���y=�\��!U�O.3�?X����6!͖�t#Ug��Q]s�`��h67�*E�A$=�~󇺨�i��$�ݑF-�yzj<��o�������
yg�Fh�����HhO����c<��*R���D��ܑZ�Śg����;DV!��ߖ!���M�����=5��	bAr8�4��CK�J�#�$��D�5�C!<�2�@�}���2'!�I��;PT��9X�|�Vp(�a�R�k����e�Ɯ�V5�؍�14�0	�Y�_m��Y �M#���Kv�TE��g��J�xޚ�\O�e�Ȑ���+� ��\Cu��t?��Ӊ�����-��uR��z�--L����d+�8�V�#	��ժ{5�s!cL��V���)U1���h����E�X]y<�Ð�PLAXy���$�5���?���*�1B'8�L�`!�X�����
B�w�ź�B���V����+wr�7d?6␕��S�JO�{�ߵJ���mZE�nY�<�ⅷ̺\�؄܈���R��7g�J�lŬ�A@m�z�k�x��q��-~;N�lZ�^Sc�Y2r���U��5C��]��+7H�!��*�#t�ߚ@:	���8��CՇ4=Sr���bG��NC�&����z�owQ��ĸ�n(�'����Io�\�g������"W	�y�¸��-]����)�#��d��]GR<�H�*��_{���'B߹܁][�6&����a*5=���GO�������)S���Iԕ�n�8Ԑv_�N����p��j�s���<�O����Qw�&�!=�tfO瓯h�tC�w�_��l���H�����Of:OrW[��W���RR�L��-[��^���\~б�����$I�t��^N�^��L��ɰT��
~� I|��;=%]�#k��:���1I���w��T��k���&��o/�1Ж K�� �%J+6�*��O;:�����{���M�o(CO��Vk�ݜ`��q�/S("\֥F:�A�|ɓ=L܆�&72ͤ��ܨ��8蠒UJ��m����(P�lu؍��5�k�M;ԥ�К�f��b�M��a ��s�?�$�V�"4*߰xkm��Vp8���:Px=����"&Ip��K�HPH����d�"��|�$vZir��{g~�VW�����ψ?US*.vGa�%�񩊑s@HZ��usY��u��������~Ăt�� ��|)x�w���o�IA���}Zׂ�������޹�;��O�����%Ed����2(�yǿ=������� ���O&�5>��h��t�O�g�ٌ����}o�1݇ˈ[�I��)T����p���$ǡ�0�����$jX3&�x��v�כO:5�(����Vں)G}��i���'�0����J�3���Pq֭�������E�����ak	�Yӹڸ���c�s�)X
�u�/21�m���1W^1� ���r96�ò��4��X�]�=VH�F�>_�#me�YV���<`S
����Q�00�/���]�}�6��dO�����f��W,�sJ7OY*y�I���Qg�WY�H������=��4)_�:J�L	�ρO�e2��q$vC}b���sF9��4�<t�P���q��r�tK^6���NĬ�-�vÅ�� y�L�X��0�M��`�fCf4����M�7���gZ2�BL��c�yc'��W�u�|�Љ<��G�0�Նc�t���<�	�'F�L��?$������+��;�
�]3ۊ�~�>[]��* � Tâ������d
��r;eu)���l����t��\���k}���ߛ��h�1���5,_��3�5�u̶�D�RL�,��SS�7�NSs�G!�G�4��
u~m�k1��hV�Ky��G�T�`g@^�j� �����Q�ޓ�(ׂ�!&s��Ѡ/���m�rsNş�%�5ybE��Nsu{��[C@�����fz���R4�5C�Q�3���=Y/�xh�����[�x��,3�� >'���ّ̟���6h�Am_��=&��?�X@������ggvK^�8M��Ǖn��`�k.}y]$&�x�6�I���>��2̙�0r�Y��Q���O��URZ�#iw�Y�Ɨ=���b��0+> 6������۵^��ys�x?wQ
��5��O���e5�u��iqd��A%d��#��	sVH�v�ذ��r�/�Lx׿���i%j	��)�ccz����XG2+E�7����hJ'��.�&V^yuaJ�+�i�$�\���̠�_.��Z�����
	��A^hE�R�H"PU/�)���� �R�De��z`��R������E����*���v?	��KL�r��Z��	��8l�L���v�H4fV+���]�S�T�vi(�E���h��h"2sI���A�Vh�5�z�=IP	��Qݾ�HY
i}��p�~�u���FPg�D����>��QFtO�7fL�ݸ�.R�/�֧�BC{,�kW���YI�e<
,����tҵ\.��U��P�s��8���d�:eC��� fr��ӳH�&H�sc�bq���N�N�ǯ���['��� �e/�6��&(R��"���$LU>�8�K� ����|�F�m����A���u��d��C@�=7m��6�2�a_&P��? �	���
 X�!h���K�?�X�F��x����J\"<�K]�7y v�G�#n��y@�=�<��V�ء�i��N�;�@K�0�[�cw�B	-s����m�G�K�aB&Y<#�#*��Ʈ�i�nO���ŵ��|ˉ q�^��H�8`@�醘kВ\��%:�:��U���V�7��|z�أ,��:4��|���'n�{\Ji���?�J���p���y�옷�Q���
�X������a����J�臍�=!a�F�f6<�O����%�_O�j��$r
��3�$�c�x^Q�l�V�*��o�_�Ɓ��N�T2ә�,��N����io!�(��V��0� 7�<ۭ��Ή�����6x����Rr!LfUi����4�6Y���w�ӕ;�B��x����Rf4�o�]~����n����,���2�l=7��Į�B��e�I�`���2N���$�޽sL������@�zr;�G] ���3�*�
���6|��+�A5��E���Ѫf� T���]_c�Q~�$��k�ߌ�̞��r�1��_,)R��'�8����}�O�o�ݔ���D��*��$˳��r�E��@������@ב�q��=+�i������:Y<�hf��eZ��Oq�|��) c�r��/ r�ۡ(j�`���w(�Y���Gs��Iv�0�W�,[y���$��DHW9�B:�����m3\E�':m�F?�͔ӺU��,�7b���J�I����E1� �r�~#
Ɏ �<	K�f~�	���m���'�OFb˿ʽ��8/Qp�0@��L2N�R���N*l}���CR�?r+�x�bԎ&�C �3rs��
Z4< �D�+x�rBv����%k�.�|��\�k�=7�{�jǩP�R�L�v�I��&���V�5&�_���٣�CS�O����+і��-u?�7��G2c]? ���t�-F�?v[̔��8n�wjh����NԖ�ѩ���ǏLz��A�&�x�T�ޤ���_G%��f���:����?��#�%(׹
�%U���;jy�\��Iߟ�K �&��Bu(HO�. ��O�"�
��>����N�9�����T8$��F���`�0ky��p�@�z�a��.<�6�=�!�;FT��h(�[�L�!���X:��.���4��F�A��J^ߞ)v�vY(�rc��H�t��/�C��7���:��>ܷu]EH�/Ȳ��A�u����� Gk����b@u��B�m�8��Ņ�|0���|:���*�`���6���0�M7�]�����87 )�0�y%7w�U��f�VR�����8�A�Lm�H���Y�^�k�����"�᧺6�Y���JN��'��+n�5Q��|a�9�Y#R��# Q'c_UT��RM� �������3�d-A�B�M����Q���!�Ydᅴ�Af��2
ɯ��0]f�����y ������r&�U��ֈz�9=Y��E�$�ǫ�6/_\J4j���v����~�m5�Z`����$#U���$^�mŒW�#4��mqn��6@k>��u���'�ֆ�qF ��DcS���(��S�����ApD�p0�s�J��s�j�벚J����d�����j信:ޕ�7�=�$:�CD��w/*ww����m��'M�mn�䀹�tC����]'�r�i�n��t�.P��e��hi��y#�.OB�Q��?�˽�hD]P���b� � x_�j�Y�mW�b4Q�h����6��$�zFǇ_��>Q3�7�ɸN��O����{ϑ�AE����6eY_T�3�m�`��rP� �J��<���y�|Y��)|�� �a���������"V�h�D=ƀF|`N�ԓ�A������Ȩ�ųu܍F��ҐE_� �׬C+
'~S��k�411L#�n8�K�QƐ����q�DTh����4��Yo+l-�-�xh&ƋDr��k}�l��"�@_�_��2�bS���nIas�$�s+�۷|n��UFw���X�1���T�#O���`T��vP�~����Z�z�X�&�S���(�-��1��PN_h�KC�`NVۂ���i*saD�l�HN	^��l*���)�^��,���1 ����t���k��qT)��t98�a@�H��PR���GV�S�yk���v�Z��/����r�g-�/�b.v���H�@��[�16�E�ó���9� BH�B��N��Ò��,	�]K��H%YY��#0�j� �����K��/YU��d��l��$�!y�'���65X�tO�j��d��v������}G���yiE�Hl�v�M�#��d�@�ޘ�a%�Hr�!L��\ �ϙ����r�뫐�~n(�pB��n�YZݙ1������S�6-K�
���,<7Ahz�aV��5Fa�fȝ������.?��Qm${�zŐ�\#9�ٔ1����)1ϥ��YA)���w�C-��|�����> y��z���F�7Z]N��Q�Oq�f[ۻ\���Y�oZ9���?��na�.�I ��]5׌��]Mz���Mx�s�T!�D��I�^�p�j8���#3�X����>�C��'����E����>+|���)�����7x]��[F9�mC�>�"s�E<����e��AE�m���"ʨ��,%~͗���T�0cx|2�Y�ϻ�cϡ�S�Mၨ��$��&vpK~f���ͱ�-J8.]�]]�zH�/�;���ٻ�:�d�o���R������ݹ	|	:AlA���Q�F�\(�e���k.�ǩ�2D�J6n�q����P&�?�vsW���*��>r��C^h�g�7�U��Ȥ'&��s[�z�_��h��N���yOG��J/[M� j;r��1��Lz�=D���쏩m��������V�mH(�J��Z��j�����)�xN3낏KJR��)
��8�U���J-�L	FA�q��wPz��W���.lJK�W��h���8j�6���� ��~䶚�46�ju� �+�
y����浕�r.��(0_y�*�_���U��F��-!Á�Y4d"�o$ŗ��J������(����5�t-ibR�����^{��]G��`�~MI�ܦ��w�+�9�$3w�����f<��v7i*aآ*��5	�.���W˷��xӫ��L��Ab״ұ�;�DJ8l��}B�+�~��M"k9�5\�w6xW��aN�gL��զ
�h�S>%iLF�=KR���Ч�
;-����o���t���o|D�k�ѵ3�M�Vm]+>��Y�)_���'c3���+V/�A�J�J���22q��;������Bα���zK������0^�8i��c��K�7�������@"<��J�ꚽƝ
��j�X�М����g�`�#Ԓ8j�UmU�P��`+xuK�VH\�n�
¶��,������1C��K۴�.�b��8m}�A.{�Mw�am�)[��b>)�>]T[�g�������^�[��� �gK�|�T1�#���d旑��Dw�~�'؇a���0���L��f��Yvk]ޘi�i�Hˌ&�<Ǥa��Çw���4z��_H���@ֲ����C��GH�j̾���+�༌�Sm1+���@k�-w���܇�g��h�2������-�n��؄����^�gϙ��ٺ�L��o��'r�,B=���w�H�S��-a�\�7�F��z&�,�$���?*��ܭ	���N��&=N[d��J��w*чZ�LT+�E�s��R��Q2X�}A>Z&F��Id���usV y�5�oC��ضմ�#t\4#�m��dIP��|D~������#��kG�4q�z�X�������׹�|DwT�k�"�d)�vx�H傧> �e��0 �5�<g�*mā(���ںW�h�����XMosf��s;ZA���x��K�~E��^l��Y�q�P`p��&"副h_����;A��d��O<wbԥ������F��nVޔ(�����5��rc:��N�y$���l�1�}s�Z�^�+�^�9v��Z7|���J��, �5/'���A4:̻zik*r����%<��šA��B��M��v�6�n�|��~Ip���ReU�����h9>x�]�*�<w!JRxI�B�t��f��ы������t�l9�0cp�r�s��9��l\�;r2r=��5���T0�MNO$<Ƃd+Cwl�����8.�:ub/��q�I%e�b�a�h�f�Pb�'�����{s�m���L���1�=��Cp��g����)&*� ^�.���2�E�MY�&j/1���De�_*��U_xt��e���w��q��ˊ5���X博�[Ǖ�ԙx���'��u�a��Qԣ�������@:����E���D�����E�e	���9t*�헕Ɍ�����j��x�J٨��8K�'4���(�w���!,��MY�*TB��bpY�W���ة^o�rv_���=�� ��|�Z\�*؇Z����Ϊ�t+Q��lgJ*�.|�xǲ��0�+��mݎ�7�0��ԍ����կ`���B���'xCά�fB���N���,3��.Vʌ
=��~$������3~����h򧝬6m�����H��5ES&�{CRL�_� (����燕C�
�)1��\�p�g�� �6ɮk�ô�����A�,�D�[��H_�?4�R�4sbh���:�A"�mТq�qp��:ǲ�*��TC<�G���^�o+*�-}�\��ǆI�wF=W��������X����PAvχ<�FSK�2�2��k}����Y�K�d���m��z�&��k�x�C�Q������p�Y��'0�K��&)�X�"F�x��9a�,(�k���4&��*&� ��وl2)a��[^Q9������v?^B��ʔ����Knt�j�=$�Me��Jc�|M}��d+{���0�@�K)�dJ@ߥ��b�u�F���q|<�����$�=у����'�qfk�N�������(+���"�G��1��� 7S�(bL��<[1��"����+%QA]#��&��`Tw���ў��`Cz�/WR��lķ�
�3�ߐ��Ȗj�H��c�A
d��V!�#�͘"#�m��a���<ԑ; SnB~��toZ]�{?��(�n*~����#颜:��O�iߓZ5�UYO�RΜ)f�(��Dok�Y������|��ubAx�R��/��n����l���I�<��|^�aX��;�"D
`[����'0M?�c	#��(�M��tJ���_�N�σ���H^���J!2�^�Z�z\g�?��*J��h������0&z=�7\Pj󹦗�|Y���iL2S�*FO�¥�P��9;�-B�n\d�Z`BF>{~��b�E�`����j��D�ְ�?�m&��}�	�5--��|v�[�%ؐ,�^�7l�!h�i���w�����Mv�B_&��� ���*�?�vA�m&$y�+�*H�N���{��K�1�`:Z$��``���w3��t.�?�!m#�^�����S�QQ p����%
u��]ft�Ą*F(�_k}�s��)������@�˲���/Ǵ}.�4�@BCq�:qe�E�\h�Þ������/���&ޢd�N��F���k{*(xrI��9��]��Kψ�7��q�D�J5�s�A1�u�d?��J] D� k"l=��g�7h��^�i_�W'=P޾���AZ��1�@���y�|�q&�q&��V��"@�sb~p���	�i�yР
��h1� ԧ��p���B��ZUA����b�E	�U6m@�7��GZ>��-?5��q�t�! X��P�T�<h�6�
Zw�(��,��|������U����s_y�vЈn�"� ��[�|�?���㳂��6��H��E�[8G�Qm�F����s�d�!|]nX�O����)���`�a�����n�*wgIp���<⦽�^)���F�S��x5�OU�P+�&T�(4r[�W9?���j�m
_lK=��v3�>$"��LA�ITLȦ�� ��`h$��x��ܽ�=���y��ǃ/�� ���G;ZG	� a��4y��f'�ĉ�
�'lR�����6=:�E�v��j5�*Z�͚g��#�^
�{%�7��q!�4k�>~K��������j���i%lp˂@����\��B�rRr��+/J�&��F�8290���s�Q &Y75�}�v��FK\ee�����	�bL...�3}��ݫc�1:O�K7�%rG��q��A�
��X2��bqm⎳G��8P��~EA����w��+�~B��R'�ܰ�&���Y,�zJ����}^�\�qB�&3'�p���o\�Z��e� �S֭mۛ���&�[��l��k]}�o��*�v�4���7��h����;
\��0N*3@B�N�^�92S�!�Mc�I��Зf�a�?����YW��W! =D�������n�R&A�8`ю��t�c�N����lC�<�C� �4ܾ�t�<�Ж�)��3��U�ܖ�9�p�W�@w��o78�9���h��� 	D���c[��cg�|��X�^}������+��YC��{���o#`�����Z���]�X��-���Z����|4L��A!�@l��>��Aҟ~eL|���`DL��8+8�p �c�L�h�ψ�[�����4[W�n�۩�F��;���a�[�r� D��+���O�$�!S�}~��'FJ~�_iM���F�����F��Q���S�1�����o[A�	�#\��H\_*���>R�z;|Wa�,�j��4�hv�&↓ 	yVq�������^eu���_$�H�����~Z�G����-���4u��/^\9?�(bѺ���S�}wB>j�].�G�<��پ�;��D��h+�q����4Ր���3�Ao�s�l��B��v��Y ��;zl_�Mq�z�# A������ޢ,>Գ7�%,�B̚�p�y�ğ�k�c��fT��͈���0�7��ƞ��i��J�!��5�'��V�X���W�NF�rX��/QGβ��ǩ��@�/�53�Ҁ j#�0q��Q�YW���l�3r���Cy��j )ͯ ����������5��kCm#GK�	�j^+ha��*��ތ�5*����6��q�߷�Ж�B��$M�	�ߘ��m��/FW�Җ~�0m�?�� � Gm���Lץ�����!��y+��o&�6J
~�Q�\��Q�G�Fv�Er����J/gV/�42[�m��Gz�Ba���`�+Ñ��~ךG�<��%�BJs���x�|��&3���K[,+�K�ƙ����왓��(�� �h��|
#*YI��ی�,��Q���E�����#y;�H��M���b�9����]��{���x
�3Q�bj����.Cj���8��+�����U��?�R�,�W|ATm�{/օ��Nu{p�7�P����]�k�1�����w~�Z%�5a�Za�%�m	rL���p����h^�� �R��^qn��j0�BS��gH_�G13�IU�O�藇u���h������m��6��Iur�^�H�l�O��ry�A1�ag��^ɯt���#��b]�k�P"������4�M8$�������-�3ͷ]�� ��&���`G`�N�j�x0C��D��:���g�u��~�C�-�o�z��#n$BӶE���)�L|zi�[%cRP�9%���@���+9�l���%'��,-���U� b�8w�Y�qѽn��z� �ܝ�[y�m�&��L�ε���i��uN�5.tđ���W�g'� 1ٛ���D��]�ŭ���Y�e�齮����/�Em��=�9D�r��/Əݑ͆���$�9�A���������k�	��l~��6������3ì��7,�Cpq:�BL�2����r������F�L��@'0�8$��.
p�)d:�O��uOE�5�s`����nyjW`B_�uir�F[�#}z��&�.k���Xj��pmh�_|{M�T�)؇,�]N&�N��<h*i���lbiS����o��O��ϩ���Y�+�cJ�qL�=�~�Z���'����Idq$�@�r�؃�|K3�;I�&ɛ��s�����~��w�"��V�T�
�d~h'Oz�eZ��(�}�c
_z�mL`:��֡os ]�����z����;p�t��D�Ճśl����N~ά�2�E����ae�"�fII�z.���@�P����93�#�jS�'��E�'���O��m��?#1��]����43,�ŧ��s��˚>�/�o@�!�vE��a�~�CL�Eά�Ǭ���	�mC�0%���c �8ǡS�W�^�~ZF�*W+F ѱ��ۓ؁�vHP���%��w�7es��zo�w3�TI��s�r��x
����'�<���I�'58�c����m�����ٝ�������l���J�ΰ��l�iq�~(�?U�RUM��q�~qH�,Φ[��#��g s䴌� ��2�Ĥx�8�Rȩ�6��+�LbK�;�%ܩ�����-6�����$�����ub�c�_����I"��(��U��:g��նD��ɳjˇ��M3��9c�ܬ� :�`�@QV.K������A���\.�|:��n;3�T�@D�ӝ B�I�hz�u�i�<m�G��xl^]��c�Stnd��M�	VV�u bbį:t'�9�hh�y�u��c$*�p���;�^^�}(�L�-��v�6���)�]>c�f�bé���:_����䮶A�B�v*����0P�B>�5O*?V�/����#KZkZ���Jv�zi١��H�%϶v�-1#Z��j�]M�B��G "�/���2�$���w7��qqў"���@����3�`��k}�c@6 ���7S�~`��(F���t��Û��)6fb.�g]+�Z&�wܠS��cMm����{���+҉2}q��l�.��Iͼ}"��Y!΄��!�BŜ"[8�I#���W�Ҿ��۟ь�n_�V�ƶ��% V������Owlu2��ϐc�K����n�.$���eD:�D"|@�����������M��G"q'L���+�n �!� ���ؼ�}}]�/ז��ÄIϢ����ݺ�_q�$��+o�a�d�J`D&iT�vp/m�?�eeކ4
ȝ�5Y'n|�j�A9���m[b�j�AoE�R�;�X�q�V18&���*�k?N�z)s�_	d�v`4۵%�"��$��ل`��"9/=Nl�]�+��8H~���Mj�< �rH�4��lլq�(�|�p8lMO="r0!�CU��6��#t���e��<�4eگ.��a�h�e�8�W�=��s�M��ٜ���2�z"��^�2<��l�a����|}�����[��{��[N�u��7�1�=�X�x!����[f8����\��*�b	M�^U�B���ٛ�~Pl�1{��h�?�d~�%�g߸����t(�T��_�m���l}v!1��K<������InD�؝x��"6��
ŭ��}����q�7�m�*�à�W����SſA�>)����b�P�! 8+B�8��G����`e�G��Ŧ'
,s���i,�
	Mw����jwd;x���AA�_��\qO�Z�?��+��Z�N�[�#W6��b�T���ϰv���ϏJ�(O�yڣۀlѰ.�Bϲ�O���K ���S�b�$����x>�H��BfL�f�y�{��+,>bvƔ�ǉ"k�5둶�8�;[�\e���H <-��Ե���]:P��Ss�����j!���t��	�]c�O��C��;f[�y����X�@cr
_
p=��l�к�Q�DG�(����Bj��eR�̈́z�]�V�������r��kŚW��i�z�N�����J�_����y�>FR�Og!�J�AG�c����i��ٮ�5�m���M4f/7�I�oxS�n �� �B�nZ�7�P ���E��|"q%0��E�S.{���3o�8�3MW&�J�&�o�gNL��.�1�L�U��)�Ѭ�?ýA�T?�Т&������荾ٛ6+����bR���Q����ĭ�ɦv�y�Ĺ0(��2imY��S�p�z��]ɍ�����2�h���h7�n�����AΈ�tVM�3i����Q�}]A��ѝ�	E}3N]�;�?^�F�0�L�[V���S��1�����=�h[J�_�����JC$F|��h3�$�Xw�c�g�E�g���q�r�V��}̫IO�~W��<n2��C���FS{	��?��9/ؓ��o��	U�	������t���S�B�IȽ>�f��W���-�[%:��	j�Y�[��c��� �
Ԍ�H�-%foF�?�|�u�A?��u�!Ð�"W�F�,�������ځ�ϖd����\��(��_/���l���6���N�\btþNԁK����P�����.x�3��$����]�R� '�ף�x~�'�� p~��?��ha�;? ��&?�]�,���1���#{k�\a��ctZs�\�0m%Կu�aD��������2�$�y�?�݀a��`0��(���)�}� �?�x�3��-�"�Wh�\:��oC���/�W3ٵJ}+k�!��^9����(���D�6����{�e�Ǘ���R�)��:i�W�+g��  	������bw�r�_���Qq�D]��L�fY2��X|R��6"Y��/�Dh>�+��GX��b�pr:��ϗf�~����r�b[r�RNO���N���a�5> �-��!�^�5�7C�9�b�������)|�+�&S!
Rx�72Pa~V�3��7>^�D �{:�2>��?P��E����4*"
*B�țl�>�zYإ
.��-�L:a�Z"�I0����O{Up��DRt�9�LR����tt�~{��\�(�j��g���s>�R�8�˛«��g�B�ԹJ%�0����>���Gx(�)�Kn�Y٪�� �O��x�^�jqVM+1e��?���#A�b��=��kOd!#�����j3[���4i�x���8���+5*o^���G!ظ�Oh���E1��w�d���\�H�o{�.�\<���
����O��n��|��߻آ	n/�\�K�H(��H.I�h���h�i��'�b�&��Y��jHk���s�V��ݵc�7�{)2�4��>�W��YE������H}�oxfN�5�%aw��B,j;����@�[�8:��}{�r���V'.έ�������\*ܽ�ቸ�C͗7l֠�im�7�c�9q����P�=�M�|ѳo�a>�1+`��zߵ��no�,_�_�A}�N]�X�����~����?E����D󄚣�~G0�g��f6����w���LIJ�~=I�6l[i�/]7������)��6XI@�Yi����� 7+@o��CN6�����)���V�-�#��bs3l�����AZ�URV�u'�Y�ʋ�2�\���'�V����mu��j e��#��v��B����$��D��8puQ�@#�y�D�����.�t'��m(���M��������p'�� ��O�5��0�����6�W���Z7�;�m��;ʙ!�1�{9�i�=Y�q<J�5T0O��L��ʸ�?�**�����ҙ��ڔ�)�(���I-,_���eC�4����6����Cb�T#��U}N�^uPTa�����J�K�g�u4O2��>т��ď	�M�o]�A)�f�V8��
x��_�z��Lr�R�49\h]�bG;d�?C���jS��R5����!a�C�R�,��j!�ow�_��e��x95^��ͽ��;H�I�_xV̱�XQV����ɖ?-�����V�ͷ,��lq'f���L��ֲ:�}{���]w�T��k �\3�Re�$>P�d��e���c����JB�Iy�w� �Q�&�E��T�H�#�nt��B�����)���i���Ur0�瀯BBK�J$ˑ���pVUt��F��n��A#��+<�V�<2!HSb�������!⳪�K�S�?������-�n|ͪ.�M�i7@�6�٬���.`B�����F75:�@�H��,�^���Z�N6��5SG&a��H���D� �˻�]�����d�k��ohAtߘ���z�Y�G�v�PUQ�jV7����ʅ.�@�t��K? ��L���V�j���������4����ݐ���<<R�=��3^��7֭���O:�m=����]W_]�M�FoJ�݋������-���`�wU��,�&	S���z�J�m鑙h�_H
wҪ�?�lpB\���/0���Ёݙ�`2��<�.B
G"��5����KR�w6��Pś�8����@&�=�
�F�y�܍&
5���>��B��|Ã;w��2%���/�X(�lwG�X�
��	���h�@Q]!�f�����G�J(�(7���Zv�����J~l�P|������"�X7�Ew�n��Y51��~�b9�������� ��$���d_�yhz�̺�8,b�46�.&�lM=]�qw�#2�Eg����p,�>��+�/��v��V��U���c��n-|��֙-tÍAZ��w�l�e��������KL�$�g����ł���mTFصp�#�^�r9LJ��R>Z�Ã���m�/�W���E�����j5p�������Lx�y��"0f��(��`��۩���I��~2289M�eY��u�AG��������a%��`�M�g�ItYJ�*�\�=�F��<2Gع�Tﱃ?� ������n�,�"W��g�݂�1�|�/V�=\�T���
������n�Bd2'\�fﰲ<H	�lvk���& G���J�5�J~�al�e�|�/����
�y���6�ER��C����x�`4��cIj�e�Х�3ie����v�8�n_v����_�����
�mQ��d���}.��o>�7Z�p-4��0��+꟧ab>w�1����6�|Ruܤ�!���o�VTϠM?D� ���ҏT6��=��*�-%��N�;Y��Y>k�ycib�gy||�Q�2s��^��dGcq�S�$Z�:=�1�V�'#��.���9�z$�V����zI9� Y��dY�`*룡3��O`;�����/!����x�B}+�0�)˞�2��F���#0m� 	P F�Z����|u�u�X݅>�[�Nb; !U2��X{�l&E��e͇{QN�[���qȉL���u�<oC���%U�o���6t��ר�m4�B�j._OJ7n�V$}�Q��Ķ%�1�Z��7߰t���w��P j/�DU[Hڨ���D^s[M�-��j۴aY;7.�Q��O�d�IY�������6��<u�m�Lq#��a�����& Y��G�,1�&�(:&܏�r5>�LDPϴ��R�Xy>h�󒑘 ���Lόy�ҵg�Y�_0�&:6�$�/�����r�EΪzj����?�.�u�&�x�Sk'�ıb�f�d3с���P�{�'���F`��\��0w��hd���9t�7�����,zg)�t7 �?��g����W����Q��� 0�˽���m���!a���R�R�~�C_S�Dߨvv�oT���3�](��6}��5+��J���ގf�  ������wH�(� ��q���WCZ��N�}(R�E>!C۝�{v�`�ŭ`8%����_8V��;5��mg���OE{=�P��j=�9�H��R�a�m���)>�Lz >n>�ƧC�l���'����B����|��B㙥I�KNb��^:���4$���_a�n=[�(OV'rn�6�����͓Q����h�L�g�a�3 ��-T:�-|W�L[,s�V���&,�Vv��]]�*/T�)�_�+�QY8h%òKy�A|ݏU���D@�A�7���n�4�h��c;'�8jc�Ë��G��L 6	.���E�֞�s����}�o<�5o��k/jӵ�x9��V��~<��o�,B6�%
��XH�IT�J��I3�#��7mԜL�h�.j�?�f���J2���nQ�X�eI`���9��d�0���#b���ߎ<�5�!�w�Ju��L.9=.�� ����j�s�>0c4���i�������tT�AQ\��*���5���0y���Bs�Ӭ���m�P�������1Qd*�k��mk����%Ӡ�QV�k�{fE*�[E	���_a^��B-���X��h^!n7�+��)�d�������+Cާp|���I'�e�eٍ�Ё�������L�>��13~jO&:�%� �w��.�wO��T�(%�n�W9牛�7�v��/Թo5�C��P�gT��(�+5g��U�4���'�MҊ���zw���0Kt<�A[�P�>d6��;���b)���	�'	��"@����s��:���~-�=UW� ԍ�����n��3^��{�s?y�C4��?���8��_1?�Ӧ-ݏ�w�i��;�K�{�	*�-hn�}^ֳD�^��I����גV��D��`c�ԕ�L�����
�FJ#�-�@���~ �����#?��ꍌ\���B�tJ�RS��g�Y3��H�eG�PPf��+AF��;��tI�f��S4�)��8��=F�&����E��٤��N}-H���D�f�9����=.�e�YDdO��^��q�D:��ȸ�Y�A[���̛P��q�r����~��U�LR��Q�Ε�{��<F�p��l��;�c��|6����pl���N 5��ĭ��}dī*v�=�-�ȴ�+i�욁����۴q_�iV��*q.�ʧCv�N�vi��	��~/�֧}�x����bFmt��
�<2|9�I�)�f�^2#}֎���S���#�"R���kԿ����t��j������8�Q�㹬mi���	ܲX��x�9�*M<i�f�jS?�{�dq�6����s�IU5���HS_Ɛ���߰}��/��]V���u��\�{s'�J����<K���=-����k�G���PC��w�_���yx_��9�\yjm+ t��U��X���B�9��pj�$5Z��A���GL��H�k�j�I�u-s��½�[0@b_���J+�3rVYH#>���	
�]?�ם(���\�0��XP�4�T��l�?y�,���t���Q�F�F�ĝ�>#�+V�D����0�4�wu<�N]��@@\��Bs�B��et����>�iA��T�y�x�;2��A{��~:a<2�m)��b@�-��Ɔ4�J2sjq	���)ϛت�k���2!�]������w��9�ҍD��8�7��t;��[�gc X�� ̸E�2>nn`ig��57�v?��\�����$�aBH U�@��*h+�Z2ai^�	J�����:?%��œdIr�t�I �S�v,�A���)�������yæ�'=	��1�#5b��@���[S�Z��d�/�'����d$�>�b� i�
�yn��t$@��l��vh�F��WM]��:��8� �n8��QbQ�|��*�1��<�H�~�o(�ja!��#G�d�汕GE��� bX,�""����~@l�Q? �'����J�x[�8�*�T���@1��л�PL��@yPf�Pw�����Wv�lB�����6w G-�z%�%��+��4�Ny&ra���lj���d����w�9����W�d�4�Ŝi!c���f�3�u�f{+ˮ��uf�ɕ<m�F�@f��r�� �J;;<���U�z4�������!*^�N^rp7��j�w�q6��t�н*����Y��lRȞ�K����rgئ��"�$�+����B�E������⋃> [�~)�0�;Њ��������4�)`�FZ�a��Zj1���_��l2���O_q'�!/j�~V>�6;gq�I??��X��!S,R����� �����piF�F��Y�q!�4ֺ��u1�S�>�xo-Q?aN���s�j��h�J����Z9�ʒ��JQ����DkN �@S����y:&�p�hW�� �SM����v�EH#��F<�܃��^>_�BP|�
��˃N��W�7�|��E�A����1��A��Ј�E%�.���@U�Q�~v�;4��CM�E���k���������f_��"M��`���Ww�s���5�=����$�Y�"y]'d8�C�u���S��O%6�0�����"y)!��]� Q�z��uEj����iLzh��ȃ��`5�M!9�&��v|�ƛ��g۬B�WR]�C��%�bC��L0yW��Z6�Rr��R:���ި�+���5(� �&����e��s�	|�N���*��
o5 �tO�z�<�s~�!�����C�6�)G���͛/�Ä�`�5�h���=���ek�\��>�^��]�W�y�Ev��������y_I��`o�<���_�0
5����e�ڑo*�P�r���au��?��S��-��Eձe'E��oz�)�.�`��=U�g��a^�.�ȕ����ߟ�5�<p�M��3L}��Mݴ���ڑ��
�����Xհ���lsk���7���� ���O�1�b���{yh�p��JKy�L��qRHD	�6&�+o��/�xk$0����ǰ�G&_�0~�4�+�lT_���6��)���[e
����ӈ�c|�!���f��&����t�̲v��G4�7@q�
����;)j�%�X��*D�5�������kZ<=�4���Ԏ�R��Ӓ~�yr�3Y;�z3���8�2�J����j�� ��>٪�W� �#�Ht�0����os���1�!�E��SH��/����
�S�SO@v���O��gD�/T]P����>���a~������-���FIww���ӳ�����#��ϼ�-��^0���a|0�d_�A�:R$(�����죵����;�i"[�)�1��&�C�S�dg$B~��	E0�L�;��0�����_^��u|����l2{Ʀ���0��Y�L�ǹO�f��=�Y�IC@��43mʋ�"0����}d�"�w�G7x\܅$�)?�T��#�:��l�_ b?΁A��ƈ��Uzo�?D�� 8i��駍wsm��V���P�Y����h�_��@/.��RQ�5ۜl�����o�x�,@��&Mi��լh�B��g���=̽Ɉ\0�ON�xb��U�j4ݱC�	f�x ��6���>�)�V�?2�׏u�ee���V�z����v������Ǭ>����ΊCVv6���$��]�o�"u9%��V���F����l�wHZ�Z��}b$)w��HP��}�Ǜ)g���۵���W���L�ƍ�c�w�!Hx�Z�pnkB����l3����fhi��y!�-3w��4���M�;��	�����,�>��
bKv`��3��QO;yѝy�U�}��
�
g�!_�ۿ*�qK5LH�t(��ٙ7j�j�^D�X⨯����4���k�������%w���y� ���,h��]�p��e�I6^z?�i������
���f�K����� !���Dn�w�a��|8�ļ�����(�?��}A����XȮ/����-���-�}8� ���bW��Lŕ�����V�t�8�ğ`�䜫�:+�N�]A��Y*�N�dwnk�4��V �����Q:21X�+�6����j�l�xQΊ��=�[��"��&�>��1��q%5	� AY�L�PC��v��m�����	q2S��'s@�%�0�DR��%�n�0?�'��TIX�x����`�ѻy�3�)��MB��e(c=,����w?���rGX��BuJ8Y&���t�ڄxڋ�Ĥ��xb�N1��,�eۇ�B|�1��Ǡ�^:�̲q���F�:A�� �ר��CÝ�b�ns��G������׍��(�@��"{����^?���E�^5u7e/_�ej�H�ڡ}U�@nKQ/9n���Zh�2֞ /����<��g��˂��v�l�<�׮�p_�;�R\*�7㣒�[=�l�a�<����󠽹��4�$�+����?�3T��aN8���5��u�����Z�ݹ�67����O���M�a�g��)<�]}�#�S�rjgd�[���d�҈�#;��;���� 7>��28@n�{ֿm�u�y������vظ��;%��Poy`���U�l�ާ$TSKV���M�p�N����B���>��EL)9���F���ӂ���;�#���⃱���z3EK�g�G����*�=ؘ6gG
�lN;�K�A�k�MP$$��@H�5l��L�@Q'_�C�By�S���P#	$�%�"�5!���RH�Gx�F+J��^������3U��j��-��|0�Q�{X�5��-�A�6��vւ	22��ɓ�x��L\���i$�c��Т�GnWE�������k�����S�:O���r�G�`[�hA�ޙ�k�O5���E��;i�P,��n�74�������xU�XN��D ��5bhi�A�
�P���,X��mjl�n]�$�g?�������QШ:��Y�m=�þ��Y�ٿ��5(?W�u��x�⼔cjѽ�HL S󂅑�c'B�(m6�;V[�׿??�8�dc�z�D�ܔ��1�|��:��1R�G-���yh���/Ų�8W����uPS��
�P�{��	#i,� �k^t��|�,�b�UZa����h��'�9��u/�e(P;'o"�m�~��r��˃4�']�L3�v�0�'&���:I������p׉�H-0��b �wl#�.BYNj�U>�#������ֳ����KZ?9���?m\�!��y(c�n�.�&x�#
��	z��!S����t�Ʊ7�R;�����;,�GzS�;s ~��=��U}�)�uˢ�����' @�R}_U�%���R�U� 4�d4U {�^:�ھoP�+ qbuY��h1-��r{S�VN����[�u��
^
���@Ӡ��V���J���-�.��j*�K 7z�R���UX�J�Ʋp��%#�.�Jם.u�$�ƿ6�� ʥ:�lYk�0ь�-�ҙ�����SK�}<A���sx9�)��m5��.�O4��s�5h�&4��6М(�m[M�؎��'�p�k�����z�!Ѩ}�ч��޾T���˓�}2��6�N~� ��0�]����42xo���s�y1[<�(�!���fӧ�N{
�&�����tqզ^����p:���}����H(-aS0dn����Q��5��Ap��˸r]N Ƚ�ϔh���1�������p.WO�,��f�����E!�����dƘ&�o�;$$,�rIM�[��2��3v�E��Ӎ��}a��V���K��۽���
�t�ƣo�O��F�P�ɛ�5��*��mxb]���EG.Xj2V��V���^�����7��T*?w�!W�$}k/%w�����
�/�u�D���u����U�d4I$'.8�u�j�����݊}�s$�-���4(6���S�+��J?��#Q��.gD���)M�燹n+��_�4���,v��H��f�!�J��]���?�Pm���ِ^�(oEQ�/�]=�K����a���Y��)���ė�@�M֘�X=�l�;��d�@��F��cQ�z/�ʄ�WD<L�҈;�`AGgE��K�'ę��6����-QܸhM:���*S:�N�:��������M"v�H��,.'�E�1�$�[ua��,]^Fdߣ>`}ʻ���:#@̛w����a%���9aЪ�������/8n�ġÓ.�q�g³O�!���x�B�(x��.�����I�3f�����F�⒛��v��lq)>�J�%�lY(�ުl�(MH� 48�r/���H ��h�*a�iHU$Tb���ivfFD�����^^O�ױ
����0���uj�Z ��D	ƂO�	�M�@H�iY�-͍�-�h�=�3��������QZ=�+�X��ɤ#��*�s�ej��4?L����`�}y�1M���+�p���/{��׍!��%�������2�I!B8�L�5vOل�]>���(k�&���S�3���o&�,�6>��n�N�ݠ���{��q/��<O�f��.�{���nh�f
깲�',��?�A{ט#����v�v -[͚Vm�؄��
�)���`��ͼ3��'��`�T��C���A���	�ʿ���M��;�22!�3��U�Gr4�-�=�y�����G<F��"/�Ŗ�.���E%�����i �Є�?m��V\�zz֛�n嚙ͩ�n���ԇ\�3nhRPF�-�,�;��X�1L�$��h�P�J/��n�5���*IR�e��cɖ�V'�0X�� �­ٱmj��r��v���X�eA�D��G���s�S3_�!+�l���������8$י�����E.�HNv�Zp0L����ݑ��5����hn���/��!!������w۩��0��\�b��.������I��bC,I��YI����ԓ����t2�!lY��b�!/�l)l6`��-�L��xH,%�q��pg�Q�_ P忺�7��.@떺C�����p|�/Mg�b�,��~��h+EKƘB��V;S�e��j���N����E�髀6B�W�!a�A���3�v�t+Ƞ^���&�|wA������Ms*����C���HRy�%���\��ސ��ۙ^��\��.��<���d�b��@?���T��Qχg�C^�Ծ�{�H��E\�gj�j�*�2Ư����/��b��<�>N���! sn�ʢOn��1���Ьb$#����,�D1��l�����z��I�8�c��u��O���m��z	iF5j� 7k��0�Q����f�'xI@��Fx!IE�J�~b�-I$v�4j�+�痲�(Z 6���7=�-	�Tn��Z��ex9��/**FeL�L>^=�h3�W��Ebo��y]�U�b(C���7�V�f~gK1C;�C}&�|w�#uZ�-�l���%�V��?@mFګ4u��M�(`j6P�hݮ���q�����4�%�X����@�꜄`�7�ej�9�U�����b�7#_Օ��
@5���./���
ܣ���U�貉��cvv�B&���5u�5�st>:/�w��2�z��W?���89t�d������&[�^�1�q;x���n�!�g���[�s����t�^����.�o�"<�]~�@�1M���v/.�#n�f�v�>r^ω��R��Wk�w�*�7�r&7�6�Z�_Fo�KB��:�pR
�]����dt�m��Doϲ�J'y��N��h���
{�T�hل���~l�g�y����Zl_}*��Z����;	�<�a&���@נG�e���dL�2K�k��,!�Ra��0P�u�?Կ�f�V��G�Kq��~I���L�K%�6_I;��/0�j�5�o)�d�d,;���kW"���Y<K�C៦Wwv�ى��O}�!�G����br��R�2��'�{D�`����J5IWFo �V����.��6T��g֨���l���aW��o�B[����<,|��S�.�2�g��{^*!$�J�Oq9M��=6��ޞ8t2�@��z��l�[�~a~�>��/z���++@��&ȗ�t���"�#������]S��"���][dir�Ō`{�3L}��=-]?C���c����0(`��|�v6xMm�k�)���umi" d&����w?�Q3�?-�ơm]}\��߾���b��������Q�1�����ws8�Tރ�~�n��@{�pU��8D�gw*)[��$�q�;�`����M�h��T�ָ�2�=$��[����^�{�O���u������`��[C穅Nłҽ�v�ў?���H��1�2y&�?Ԧ�F}�|G!1�Zg�8��e:1�`ۗ��S�-�qo��C�>�-s��@���d��N[X�ׯ���\�n��fkG}�����l��#0�Fn-�����Ns*H�sBŘ�"Pʵ�I/��s.¡�� v,�iv!��?1��7�W�Ͽ����IT���$:�eW7@���K���=Z	]	)�_w]cʤ;�1�!Iu���|��J�S��������GV���ཻ"2Eگ�ꇕxe�pЀ�oI��xʊ��"AY��%�G{|c�ؚ߼�{�[Do`�|Yk��MĶ~4�ȹ�:<����!
�
+,|�$�sa���-��"[�5O>�8JeQ��@Η����t�M��@�xzꡍ��/4K��Y�%����,y��т��uc�;��Hܦ�� p�h����	�?��ظx��B��D��j�a[5i����+]Ip�K��hǶ��n�(;f� ����gRaSLv"��w������˯w��'��|�덕0s��E��cMl|��if����0"~s�Gk�����y�4Ń��G`P=�F޴R�^���s�2�����_��"C�S��F@��c���
61-���"��N�n�3�Ӎ7x��U����^x���#���e�6)�S�[�B����,��_~T��qp�@|V�z�a*l�|BO�r�;��c�N�K�|�	B8�E��k�|�m����Ri�7�����v��.��9��Hd�~[�[�.����c��@��A����7�������F�ь�obbov}n�3��v%.�柪�zJB/L|�-��E�����BB��iU�w��V`p~���V�B �EP�Sh+�L���X�FQ�P�A�|Gf�K��8��+�~q�G�5�k���d���f����+���>��ђ�z`钪%F0��,�+ĝ<56���)tyD ��T�2�x��]>�6?1	�zٴX[��~��v���J���A�P���գ�ѝk����R��)0F)6&M���4�j.L��^�j�yM��M*�D�� b�-EVr[-Fm;8|�<��#�'}���/�&�6��C����eIs��f �����Zu�y�(rhR@�{��͠��[c�N����8\����3�bN��O_�(�S�h+/Xi�`l��}�.i�:����%�z��oxZ��*�����>��TV�JÖ�F-g����d�c��yV��)*uҊl�Q�
Я���0�O�Oh���FV!G��w)T���B���ִ����VqPf Y/'l#��Ij�z��!��d�6��^���"uf��> �p�mD������ �/�d
XV˖��Iᐛ2�)�Z��
Gѥ����jQGh!ñ��z>4�%�Xc�qŘ'Y��q0SCϜ ��~�ryA^Y��v�p�t�da�ڎu�{VG"��΢ �Kk�Ԓs��A�����1�D��D�iI�R�:I��K�h�9��yX3�w��\3�U0� ꠽��CI�qd~��J!��A=�A��ҹ5�{��,�5[�v�}GH���
��C��Q��S*9Fn(t�����Sԍ6��Lג@s=�Ê�tQZ O�b�馋`�:g�����8n�����UMl�c�!�R�`�����mQ*u?��-����~\̾��F�}9�`HP}8}����~
`��Bvqc�7�̀��$���I+��;B0)�3c]�R9/!:���z����m��Cׁ		�~_	dI�G�GzX�v��
�v���F����0�%��K�P،����2Ptۖ���fS�:����2ܰ�����m�S�����Lw0�
��O#=>j�~��H? ��F�	$�/	X��gYx���ӉtO�{2�G�d�/��^�tΣ�(8�j���@��*��F��X�ʐY�
*VM�ü�j(�qƙ5�fu�u�st�g�ŖBH�grt��O<�^$��a��������z�R���o�3�,q'��%ШPD�c�!J�|~�\.XMVw�"�r40Q}/����C�Ж��X�Nt�frIH*�:�V���~t�C�H�Ų4!����{*I��Gg���V���z��BW6���3��`$���7�{R�`��U��{mh�����T�j�%/Vc��٘u|��i��O7^��	o��%ܲ�Α`ѹE��oEX*�=Z�f�b]�������7�g��w�z���X�*��*0�VX�Q�|���i8[�I�y��[% ��]���?��3�k�]���M܎q�2^A�(Ǒ�8&��6���a�^?��6��S��]�R�@�|L
�j����ӣ��1���ֶ<0aå�r;�R[�u6��o����G��a1�F�p�Xu�a�i���O���ǧ����a���I)�a*J۱ϳ�1Ҏ���f�T�c3IB��W����f\	�}��'�c�(�]e�v�y0���H�-?k&���GT�s2�U*�]#w�����An�R<ȩT=R��3-59�����uz��N�P��	4�-�H��B�;)�oГ���� �m�N>��?��d+��=�_�W{��A�;��YX!��`��}r�m�N�B����Z��9Y(�4�1�Wb1�В3/Y阱_M��&��«�z�3�}��Ԍ�R���cnu�C�� G�	��,�?ª����G��:����3mv����;�i��-JN;�N5�����6(���
�m��l���@ț�eH��B�m>ŋ�˽ќb�1��.�n!ޢ�9��-"2�k�Y �X�U����hĄ)�`���/2��{n�iU�q~����k ��.T�Ag1��R�d�0C7��c/�ۋ��.Ǹ���mβ���|��g��m1�u�:�W�x��Fa���B/nbI4DlG�h�r3�i¨372���``WX�QGZ��;BT���(��F-����>;��WJ�ZgƼ��V���@�J,r>�7B����l]Vj���X�+���3w*A`r�߶�����*�MR�?�p�σd��&�bT�k}Y��T� n�*�V(�$K�4��x*^+a�Wͣ�h�R��lpa�xS��5�a��� ��k�U�ܬ)�w*�+�Ifno�a�WA��0^�hW ��|��_N5�P<������>��R�w	�6�d�F*JlҹMH]�y�"�����l^伿�������V:/�r"չ,E��C7&�����Q��k6i{�3��a�(�ZN��-�����L�����,i�Xل덬���5�n<N��_������<+�&�n�)���0 ����X�����T���`9���j�<2ݽ�'����P�5����GCź0�n�UY�~!`�0>�c,�F��Uӓ��8i�	e�:B���N�r�LfD�+ީ�?vk�~\��>���D��;���d�b� yؒa��@�Jf��5XQNKW�$ţ�2#E��e��pֈ����I��ݭ��3Iay9�X@Q4~���V��N����;���b\#��kG�6���X_��·Cz[�A_�d��VS�bq"�����<�o�@)�1��k
����H�DO3 2T��9�	�N.�uU�Y�7��]cs�%vP"� ����V����@:��B#w�c��k/uG���w�󆌾J���./9�{�8Q�d�9A�XQ� �(z��_��V=SZ�b0sT�R�o�E�"O/��螲 T}�p<�׿/+XQ��	���DްꋕaP|���f���U�4ڲݧ�z[�G��I-���NV�W�$S��oh<���G�^h�n�{�@�g,�P5;L��-D7��$XAۼ}� �����^cͧ��)�����]��u�)YgHH�B�[B8�,d%^��F�@��ͅtj��U�eĲ5��gr�g+�4������baF�CF�:K����J�cRa��ߚ��&k{��*pv|n�bl$�(!�}�����s�X�H��� զ��[�E�9�8<����K�S&M���4?�@�s��-�V�d�
����6�Y��BD/��Z�{�}-��K���&�^ki<��L� :�Z~�l�ֻn�zr��B�Q-�Ji�Ϋ҇?V����HX؛����X����%	K�ν{�"F���D�} 5��m䊗�W!���nƇH��sy؄�\R��+������i��}h�>����1X�.�%ӽ�n�nI��S��G'�j�.�g�M�.��1����Osr��$^�\�t����5nPM�����=y��[h_K�:!�8�3o�ܿ{�^�[rmN�Ŕ��T{Z�9c8:U��Z��时��.0��n�7������ixY�����L#�IZ�߬oE��A����cD������ؤWR�[7>pHM:��3& c����P�%8p,[6ܪ�0Ğ�uӥ�"����,������E#sZ�u�B�W���q`d�޾�N�T��B0݁�uS��c��F�t���[L�7*��IX<6�ꤴG�Ya�
d*��&��%�tK���,�{�����B0����cP�t��m�vƭ6����ƣ�����}Ku Ю[�r�a1��>��{�7��X�Q(���������r��\�'�(�e�Mq^��a�$�PeZ�i9Ua�G���،��~��4��B�.��
I�Xϒ�;6#��!��v7�� ��D4g���Ɣ��P����sO��y���Н�L�O-50Δ$��������lN,����g���Xt�M?ꞟ�-�����F�뀓�ȟy���ADHw3B��G�)�A�'X���!�3����愗K�����	Q�2ы�\��vz��a��ư��s�J�2R�)�چ���ގ��;�z�k;��ѭH�Q��b�G�Jm�@J�vi��'d�#@�p�n�^[敤gЊ��a�;1=��b�WRQA��g�]��}Nt&q�כ�G�SNndzAm/&�Ŕ�B	��e���oJ�נ��o��Mӳ��(���d%#������/��o�)��ۈU�P�aα��^&��^\_41��gG���Y$C�B�^'�|�Q��?v:W��{�p�X
E�����m���F�� �2�v�`r�cT
� m�:���l�D+m�}'<��o��F%���t�T��ЯR5���5�z�0�J�f����,�G�� ��Y�����r�!��!�e��}���,G��&�����R;�ե��|U�� �8`��˄�Y[�&�2;h8�Fr0@.�4[u�-=�K{q�]h�J0�z'CO{���c-����D��GZ�ߡ{'��������<���"��K] �ԣ@�Rp�*��#ؤ�.�����GŒ���UC�ġ�:��y`@�XYT����@�9%�p��=/Ho4�x�1�y�n�z�����Q~��$��#�U�iE��#�kT?ܟ�� W�mS1�b?�bS��T��b�I������z�'Å�!_�ٽ��vq�p���&�Jn%���ӷ|w]�
2ѳt�[ɅO������Ry����y\��r��x�̣�R  +T-�E��$��`���n��g;�2���fV������^�3��Xe��Wx�v��Aͽ!~���Q3j�ߠ�6�Q��Wb3��s��� �
��+����@5��T�T��X�ce��WJy�h�������l�����L}�|(�@}��g��,>̍	U�~����s���F�9�0Z�{J?��V+T'I����z��V�LS����~���:�4w�檲]g�e%~S2����Ƿ�Eee�t��	�d?���||�w�:��*⡹�D��޺K+.�����m�t�����PE�I|:�ʴ;3�#�aD�W�n{r�T�|�[�4��|��y��/F��/�.����{Mc���a��-���?��E�z����r�U2t��ʗ���
[*�=��@C_�I�D����3�r��\�K�P튦��p�|#�aRT����R�զ�C�If�W�_�_�"�M�ѩm94��>��㟤	�d�*��i��L�1��,�H�͢��M��p���V����*�#DN��_wAA*`�\��P���q/C�/u���ܰ��[��h j�״Yg�!���F�5��b����Ͱ�`�9N��g���`��cX@��Bb���4�O�ޓ��P���}���jg��O-H�8�����q�iڤL7n���SZYV#I\�B�zVן����,�[$T��_L<�o�W�D�{�Aw��ti�h?�z��5M�9��k��A�^���T��<1��<�T!�1�	r�l[���WQ�ޟ^T�u�!`?��m!t�y�Cߥ>
~������-
�=����V�1�Uܻ�E5Yb�"bf���3�R������<��~��+f�R��DW��z��f�#U��M.�;5��7U)+do�Z�(8��7=�D>��
!g���w��*���T�}-���Sɟ��~�x|g�45��}U�Q���d���֐�"nW��.����M�ҟsb��߶�#�S���Oط׹��й
0Ί�P �������1@M,�K�	9:��J�"��g<2W���R��P���_��FG��KKt����gxß)�4���)
��`Z;�r�q�%��x?fw?��,�$p�(��y_�\x�~[��UL��=Q+�(k[��-#j='���՛<(eU2�M^��Y��BP����S�$�C>��ԯ�Q��A�G;3����=��2���z���`��]�
t��[J2)	�J'����SA�V��ǅR�9� n�)4g��⚡
U���q��%��v �T��!�zߩ����7���W�3͸v�4[P���if��/SK{.y��:#���ܚN��|`:�E����=���'6<9�Yp2�\���>q>n��N(���:'��𞼊�M�T0d�d#�e�"�;CQixRsSA'���%*OG��%��J[�jBnO���4�P�'{�@����o��<A,���sFIU����}u�(8"���P���z8Sf��dv���w�25���VŃ���0�%)�TM�Z|�Dª�ٵ���s4�RB)�g��:Ԙ��ҁ����n�c��ک��I��p�΄WMzѵ	����%��1��^uj9��y�h�#�1N���,�]�ܐ���*_{�)o@P>}<qf��R33�A�1�14��	�ۗ�O�W��K��P�����^����*F�Ɂ͵���N�:���/n��Spr�Z�iu�3��]��D\�K�l��9q��|�e:X?������t�(X�_i=5��-�'��T�s�Yb�'��!g���n��YK �\���"�O� �p�xī+�`��_Fb�ܞ꽀M�H:��|U�����`z������Wc��[�Y�6�вNeD�5�Hb�Vp�=nVy~�zݑ햺D ������9��d���WfŎ_H4Vd��E����`ů��la݋��:��W�ag�|v��[��Z�H�9mH
��!Y��W�UUUi��wUҶ�xρ�O6!�k������}�&��/f"OHAw��?N�64�0V���#-r�������˼F/��A�KW=��)O��jC��wx��i��L�ӟ��rDn�瑼xj'ݺ���x�Q�Fh�e��&?2MO0`V�v�e�3+�����|�U��$}�(�K�r��\�_9�E+��;�D�n�"��t5LL��AI���@j���;���|���1[v���%��E���/����>���"6G-�.�G�A���0B��d�� m�>}W-+�h��m��5 �E؈=?�>��:}wYk�����N`��蠝��qs���۸Xzs��?���%ҵ��R���,���
��QrR*��y��|t�R&)_��[Te��P��u��:0.�.Y��b40wSw'���>�'��ߐ��2�g?�̓�$ҁܑx�f�%�@��� ��_)�'�sB���n''/pPymٍr8p��t���e>�N<�[��5N�uA!x�D8H����S�����|�L�� u�P�l���H��0�Hܑ�@���zq3�R}nt)$N6ꯔ!�͋�{ׅ��h����������ːSU�N�-�̎��)a��x���x�>�S,i�SÄ×�'�kg�³�ვ��5}��c���j�0�ǜW����?S�>f?���u/
���<m6�̱�
� ���yQ���\^��u�}���3@���f�����|����Xj��h��z��mI�#Gņ9��r}B/��Z��iI6MR7���S�Š�~��6�~�FI�4�����]v}Pv5���JgL�T�� ��om-+q�)�|1�t�TҚ# EPʙ�`�JV�A�r����H��J����5j<��0� ��x�T>i�?.C������+�Z�o:�jt��w4[BhO�Ts)�?���R2�i4f�����m�k�&%���ke��B���ۄ�H�ҭ.#��M^3Q
�9@��뚭d2�Vvl�H�=�h��m~����`���'� �#m� [��O�崉���(���.#<ذF�nr���f���Vw�7��<*GO�a��\�$o�+�5�|�%�6�����1=��K�_�%e8p/a{f��5r����/<�(@y�1T}��	'񆶽:P�oi�-�w��I
B2l3�H��q���vx�[�OE#�D�i_6����b]�3eN�_Bp`��6�/3�s?��9�?�xۑRU��Ӝ b���]E��[��A�hci>���!��P�vLE��P�������ٔN� �p'�(lL,���.�pK��7D�C琥I���{�)��]��q��������h�����k�Q�K�W@Y�E��րB��2�#�UG�I-�����@l���1�(s���Q,���L�S� (F��++��8�Bۮ�������ߎ��5�+{%�fWo��:#�t�f��IG����`2wh]���1�2�����K��NS1��K�lg�3�;������|�dX�mx?���,�&�3s����8i�z������\�B�Q�U�Gk,d����ߟ��ʄ�)�� ؑ��Q]�L|��oy�~�.`�i�s�O_!�܊�)z����>���M4���?��j�ߙE`9�!vR,�(��'��������,�����J�J�I]hX[*�U`{pw,��^��* F
�@^[���8�0B��>����Nܓpm1�i"�t���F
!ʸ��~��K�}�Nn�6q�.�|xp}����&��|�0�vV�r���Jh��V���!�>�v��I���C���f^���c���j�	��kF��8TC<_���^.�R~v�b��I�͘��ڽ^�N����Uc��;�!�l���5�}��=�Cr7��@�]��{F7�]���Rd�q�ra`��jN�� &uIZ0| �k����៥���װmoЁl[��e��)�vO�#6~U:����H-���
?�osc�&�,��"���(<�Zf_�,��ru.�ӱW���=�-]�*���r�t�CbIt�g+�.��o��{�Lfl7���e�̆��k��ڳ��$R���V`�ۿ�&,t\�x�O�3��w�-ٵ�ؓ��S�{�^��}L�W'Wm��o] t�t��`�Co�cުT�����A�	�$�R%���l��p��c�.�ۛ��z�d��ˉ�`Ku�D���7��U �R��@��=ڬ����>#k!�>Lz˝ܾM��1.7R���1��L��U�)n-_�����s�,��GM�[�)9�9��'�&�
[�Ǜ;�,iÄ�w�4��~4�d��j�e������b���������d���+�;J��N[����Y��D�p�P.�=�(��� �s#���R'�S�yw��\�N�7�}t=��r7��J�4�=,yY�������i�`2x9(�w����{]��<_���|u���r~`�Ú���OG���D��K�,�mX*
��'�yj���?�Exhr�/9���œf�Xɂ_�`M�*�1"�;(�$䢟�Ժ����3K��*��k�~MħM;B��,������и����S.��M� ��B��5B��KP�ƭ��.g����фEۚaC |��ј�/��<���4������Ie��w@k�ۃ,�$��R��ؐ��#��z��.hi��� �f�2(�q I�o4aB�Ǉ9"��Pj��#��}����p�q��M�k�g�D�I��^���0��2�ȓ&����҂,X�\PQ|�M?�YaZ'�kU�'Uy�Z�|�X�qOPg";��<R}�P<�*y{�^�h�tLT��|��B��q��A��qA=v��γ9�)���H?�0g��,Z@"�G-���z��N�Jïmp�WqA1V����!rY>q����j��Y�d"S%�`��E2��|?��{@3����2x���qhY�e��'�X��{��?�릢]����3=���E!Gt�(���Q�Rƕ ���Z��{�JT�H������*�L��������~ox3,��9��&��|�֍8�0r?�TV���ZzO��G;�U�eg\wD�Vp���@�׌8P}g1G������E6=��Kަ?`��,1�I��� ���Q;��0:4<��9A[����Ձ葀�4���"ow��i����s�OH���t�g������ł�L��N ��Dkh2���z�7�D]��2#��]\㎷so̓��[_3W�,�ܗmRh�/�@�s�lc\D]�_�(j�3ݫ7]F���\�0!v�`z�)��o�
+'�&�ްf���&8țFS��F��?���r���c!E�bA&ǉ�X�&*�Z��M<���ݿ�q�jIG��,���'	���o��b�#C.��f �Yrz4g��FQ��%'Ӥ��[�����^�^%{8�8�壄����R��G�Ϻ>����F�`^��_�ʎ��$l���zO��>��x�%�~��q����ah6ܲ�F���.!���<��ra��x�X.X�jj�c��4�y���:�}	�$�W�I�P��!� =�s8�|�:��3�Q�����Xzw������D�?��G%����mS�`B,ӶK�8�"7? `����GM�:c�l`�A\�:h��e�F`���/5X-���[�~���3qb;nO�P,?nF�}��g*�h�I���<}��d�]�Qܱ��&�?HZ)7u{�����/-A�"�WJ�g�1sbV4�Qd������q}cXL�>qC����F�"	)n��]_<ѫ�D���@OE��(�����%�,��n�jK��'�r+ AC���֤�H��}*{�w$��{���"�+.S�� ��h3��Y��C�Q����G	�[l	;����l�PֹqOW��{�΋P6�nf�%Ad�Mdvfc�����g����U�d�Ŀh���Tьf�kv��a���ǉ�f�{J������uy��f>��-�J"�Va�Q#.f��#O ���<{�� �K��^k\v\⸡�R�Ԗ7���,k���.3ȧ�I��卣b��'(5�����1{8�h��l4��%�_�A�����}�}Qi�[i8w*���������c7Y���	L��]�_��2>��c��H2ú�-W&�_H�-�լxkkYT	Wy�S,L�$ ���T){�Bu�δ����p)vvC7�����ʉO�6���/�T7PD-������f�تVt��_*�&����[�6����Kx�Ŏ�RB�r]w'�'Ntg���F�2Կ��)�J�1�ѓ�A�Pݔxp���ٴ	��{�Y�]$�|K�=����u^� {��:��ƏV�����r�I{����M~��[0�x��Z�V#aF6m��fՠm��.��|[5�7%���y��F�W�H>��W�Y�G( �P2ħEa�	p�z��/8l�y���1B?�Z�W"h;�v4]����\���/EJȁ�4?4�6��e>���x��X\��n��˜�ȸ��S#+K(5q�ѻkHQ���^Z>��F�+찯v�:���q�T�c�6�`F��ɗKR�ȣ��f��1�L��c��M�q^Uk�?��YE&t8�@��]�Fì�K,]���镧��]}:�/w�%�9���
w� 2�{��l�]����o�u��:ovKH /�
Ʋ�x�q̣d?�鞎[���j���A HD�	�6�)O;D{��+v��W3x�3�͘�1cUv%L6c��ӏ_R���PVp-oj��w5	��1�;Z_�o�pǒ�w"I�]ͧge��y�[V�̷*�I{���a:PV�r�]<���Vp�e��W�E���T>@7�c�{�08.�-����xjR��91J8���Z�̹��7a
dn�?0C�&�P.��.��t��c8��K��<33�f	e,�+�~�d��ͽz����n�M�PA{�Eqi�o;U���I��>���Qc��+��'���{�;䫎����bN�6�G��#tyzbP��ޛ8b��t|OXV� ��|�4�**��C�<{�NQ���+�t��R�-�k�&1�����=�p9�h����M���0���*(���|����f��j��c���'��q��<,y���j!0��$$dە��'���vR2
jopLl��@ɾ�
_�G<3<�\�k�U+ɦ\�g���l{�&���j�"�����9�2/>j��0�wXR�G �5:�xK�_i��ޜ��A�I�N%M���q<_~<�N�{���0S��ЮJ�z�Om8�o9����V,��u4�&"|d�R#�X�>�<O�	���E�3����P���̩DF�BQ��_.�s+�yPޗ�!�aYr�+ �����`��. qK:�<&�ӹ��g�:�L�Z�oㅤum�a���l#u�5�Q?�.yI���o���z�:�IBb'��\:~Fշ�(�e/�Ga�U�I]��1�6��ſC��_@�kk��d^~��3u'�9�u�`��{����'��8�Ģ����@�$0N�"��Bvs!��<=���=������c��)0��$�{�`�J��n�nIѨ���d��2���&z��Np8q��9�Pl7��ț*5�Bjx$�׉ף"��������s��o���+�\j'�7����Ұ)~;�'��3�Ȝ�_}�ۻ?���� T�,�Z�m"�y'��)�r-Sse��'�Gj
�.�$~�z��.5/���CdA=�ײ�U�+w����)vƴz���&3���D�q����?pJ�lk(˻5�N�-�f"��ٍ������'ZaT�*l��{"�M]R�ewd<l��qt��]�{�2�Ϗ�x-{FH��ݤ����[�=�7J4;Bb?��&���Z��s.���-Kۑ�D��XЌ7K�b�g\��_B3�8'0��	�zc|�f"�\���x�bJ_���}\���O��ɗ�#��)٪w�є�:��񕰆ܧ�	'o�=ωωB�ǁ�p�F����8�>�� h<����q5�&�x&���)��mOM�~�OsT<���x���k�^�Vzn<o�'c)<��7���/^xMX�Zo����1�P_sb���np�@��?ംw�,Tk2���
E`���1
&t;�|���o4�9�j�F���3��Eo�xl����wS�' ��lw��G����c08�ވ�#���\�"��)���T�n�]�><RU�A96�Z�Ùm��-�|�[��\��0�Ʈ{+��=q�Y�6;���Z���o+@V�N-H���ה���;.�s�#��'���yOz&�e����8N�`���������.�s���Y�)�yL�_����𒢪�T�:qN6�y�0/�d��L��4���:�c��Mhi�	 �c���hȵ<�Q���E�\(�tդ�&�[z�V�!0��+I��E�k��M�xqr� k��C?ц�>_}q�#��␋����L�D���� ��9�g��O�ʪ���9D>H�R)Z#�PN�㙾���ٖe�t��G�|�FI��Gs�b`���b/(��a4��Z�>��jy���̔$Tu�j�<��>k�z�,#V:�[�P���K�/�q�¼u�D��ix�&�N���-@'�B'�,��a��3���/I-��P�#D�5z�N�P�Xt]_lÒ�8,���-
����)�5TA�QEw�qG�"�E���n|1P�xȃ_�-y;�dqG7�HA#����䏔��<�V��,E=:�s&����,���[�/�\��������M){c	������3��ȡ�Z��W���@�'���yV�i(�F�9cd���4 G�g���1����@y����L�"�Bs�4뷩y���07�p�!n��E5�U��E�G�Z	ч�;��/����qХF���6Br�G ��V��/�V�C��o�qtx���z���)n"=�Ӫ�+�QV�\��,*D�~���ݜR,��g%3>$;�Bܳ�2M^���
]��<Y�if'�99��	
O`�]�I��-+��Vv%m:L�I@|-t�+u�>�x��tڌTh�	�meO^
��>
A؉Si�����ͬ��F�Dٶ���t�ڑ��wBĴ�K�/PD��kП��Ba�.�n{ޔ��P�o_uܣ���գ�֢�b��e󿒽M��)�<�͔�Z[u�'8����g�z�i}����̇)1R��J�*>�N�R2ܧ�0:�BdA���B�C�lcfo/�l��ڥի(����y��y	�rE�E�U:��%~�\�x�|��3�1xg�'AǮ{�:���mH�|p�9�I�*�
�#H^�O	O/�h#]����I됍�@M�xr��e��#�7*ܬh2o�MS��%���ЋD�8��T��;�`}�_�77����Y�#�6Q"�,��G����}6f�|a\�e񇈱e�;^�؇��y���2.v�6r�aؖd��n�^�\�T<f��G� 2��~�b�����}�O��ï�L���ف¨��mbQ����N7p񀥄�+���#j��q���ě!Ӆ��o��H��HepZ" ��	���@��N� Xt����Ǿ��%���,�:o��3���&��u/�ߏ�'�-�����ѱ��-W���+cWyOR�Q�UD@a��mRT�o�h�[w ԩ��~2�jKd�$�S�e:|Z�n[��0��e�w��@�y��7�_�� X��x�?>�'Ǩ����T���������Ϸ=��N��
��qz~��jWFqqV�>�_9���Z\ԬH:*	�V�Wg�z\+xU��:ٟv_��(t���:�)�j���W�C3���%!�	{��<�l��g+t&r�����+�?Bd<�螊B��ʵ	�h{D�,�2)�cѱ��u��(�:۪����y�C��6�¬{����(;�{"U8%b�%U]�N�ty�tN������oWD\�:kG��Gu��}�Đ\����n2r��ތ��C",4B,q�e��^��	��md��tsv�}�\qH��w"�<����֔� ��d��ڳh򄖨5	�a��`l���e�֥XX����q�X|T07w7<8k�-<�:+�Hwx&�Ad	'�sQﳊD�	��ӥ���vF�����.�2�\�:=�Y�%
R��I8n[�o����X�H5�3�@6�X���4�*a9�x�k��+DW����o[��u���H�����J�X��[���R��	g���#wu��G�d��Uf��	�}����4YT6�
�K(}.�(t�g�m�3�uU"�v`����c�y�9s2����lS��8�3z׏�K����P�XV!��@�Q�@}-���+�P��ﴐ��j˘9�[F6o��R/��כ���xF�>�| E�8��&�f�k�5T��3 U:�����������ʴr����tRY� ���j���U�R����6#�-Q?��Tg��J��y�wA��<D����Y���c@�	?C�[4t��np�Sw|;�2w��٤8n��?�)��;��P�R��Ϡ����[5
��ac��E6LBтo����r�Dћ��-R��ms��m���Sf��v M�	0} �Aުfk�GO�q9����\��w|x�����!���>'�% ɚiK��AnEP��.$A��9��?�O�df!om%�.g����GH]�&�hm�!ǚ�R(�.%y*�:`���xv����G�\���?l�>�.!�^~Q�����M�	���8���ΰd{��=#��pw��1Yvf��$x�������kB:�_���F?�y�̼(�ZW�%瘲��G|eM�q��@f �J;s��1u�y�I^4+Aۚ��r4�:��@���9i?�v���.����I�\�����x�G��Κ�&��^X;%���̿n����}��D%k}����F�<I�=J\Ҟ'̔B��5g^���$�pl�9`~6�1J��Hΐ�|T��.�����t�앨�� �����)K�Gρ�û��%Y���f>(O+���0�-���a2О�ʽ)j���%m-Tx����m�#�T�sm��/���tm��uM(�T�bl�Q��fB
Cui�j�9¥��T#�������δ�H�vɦ��ǜ��<�؜(�<�05�f��rAz�g~�Q�C�!�j�o�l���É�u��${�/��E�p6���8�Ηi��ZT��X��HN�j&�Ц�l��=�@n�=j�!���|�c�hT�~ܽq�'��ZJ�_w;���z�XzX�j�^���a���<�^������wI$�;�l�4H#g���&���^��uR6����!�f���k�f�����׃����������ـܖŻ�e*NcS��3@$sQ�V��}���X�*�u��g���ʊ�z1C�\��e�bdMz�ޚ]7��h�Ŀ�4W��6�xhe��1S�q�O/��k.�~��Y��7�9�:����#$��F)"��3��9/���o
���խ*Z��ރs"k�Wc�m��њd�m�H�(Up��į��!ӛ��?g����.�t6�j�Q��;!�3ve����}�h��^��W�B�v��e�iv^�N��QB�xh��N=zy3E��/�`��������Wc�u�|��\�F|��l���������rȎ���,�zd]3�ˌ+ڐ~�,{����H�Ⰻ�D��;}����H��sbܭ�ǆ���0�A���ilmʲtU�f��(�c�'%�؆�'W��rp{�0nV����L������ZbK]�h����b���{@V�Ϲ���<E5lP�i�Ѷ1 ��%&���>�)|�/p�$�a,��?�&�+����#;Dy�OB�̀��#�c�?�F6pa(l��0/������-���Կ���\��7��J�:�7�u����aw�'<�qԘ����H���._���1�Ճ����a�ߗ��c}>�\�r� �8�J��`]��'4h���������E3a �KH�J�TpOP��K�ԕ���e�0��Z�EP�Wk��cn�<� :]��.y@K!���7(a��DȐ�Km���Ƹ��� \5zJW�Yjr2Ɓ��H���dJ�eaG�Z_l	5�kw6��"��6x�U�)��� �'�"��VB�	Pz����9$}��_ߣ�lU��d���Յ�)qo�.�fLXh�&qZ�7��)gߢ�+?c^w D^��ztW(g��q��T�r���h�*zQnږc$7�� �٘��7n���yCQ�2M����.*��bV��f%c���7/����fj��_�<�ES���_�?�^�T�|c���W�wǔ(64��ͨ�_��<�,�p�l��5�P���F���z���n���x����7����d�a=�/I���<
��;K�I������A��u"Ͽ�Ҍ�W.#2�rG�:T����ULװ�j��5��
�nf�R$�m0ׁBfP�绔7����R<�Ը~��&��K>��^�: #��ml���R�:���v{��
7y�Q�8G���I=Z�E>b����ξ�1:]��^�"�۹����|�f��y��1
nިO��J��?�0W~���O"׈�ʡ,��,LI��D4����;�u s_��O�`��e�<���mb���w�U�<%��k.1�+��d.��Vƿ��kXE���ڶ3��Q%Ro�F�փM���'��,:fq��eqæc%�������a�\ڙT�=<Np��*���7��V M����Ac��AiW�荑�����x��dV!X�#t$��S���c�A�T�3�kfZ�&�&j�r�J��>0���N��pCw�r;"���Ң鑎;��y8��RYM:>_����Q��(������6��G�SD��m�^��V�
�34+
�	�LIp)*B�I�(ɴ�w�+à����÷8	@����dV���[˫�!G�_HϚDi.�cŮ�1��i�TbC�(�hq��3���`�W�+��{��@6�O�P�'@�fR���)wQ��9J� $jV��2�������"~٧�T���3Nߧu�n{TV�bpab�?ݵFB�ͧq�Ɋ��y1c�Mk͓������ӑ�fd�a�� m3R'd)M�	#����H��$G��HH_ٲ��'M�rlY�FYwj:�s�����*A�#�S�#�6<���5�&���Q=
[3M;A_e��6k���4��wk���o�� 72��B�3�,\_��?,������ePh�JLq�Xy[9A��<'t(��D�$�%���%D&����܉L3�����Ư�"i��7�,|�@�=w���2��L+᪎̓�*�_f�Syנ����(J���"r�L(P UQ$O�ş�u��	9c�{�H�w�/0��SI���֘g��a��A�T1�^���;hչ>�kPW����|��Pl��GtF��h8^�Eˈ�{A����]�<����UV�o�]o�[�f:>5�Gs!q�����P5�ȥ'���,HZY��Z�>x�d��0�,��6�Sc��$[T��}̚��;T�{�6] �uOĆ������~��G��MM�N�O0A^�����3:򥍋7������tE�;s��Wa���Z�n5���ӑ��R�z1BQp�:�/C���x����������0s����4>)�z+��M��:S������vl�~^��F��K�"ѷ�c[�MG��eA���\#��?�a����P�)z0%�$ƒRϷG�A��
����5�����?w�sK�hgا)��L�#�麨��xJ+m�0w�>�#Ŭ�K�U��Y�J?"4'v6n�E�]��O5��$�b?���qi�T�U{�_��J����D�z�3]\��F8#n3UK;�&z���o��UB�d�����e�5;2�޴0����٘e��)�^�]��x��ë��6*�E��&�wSL^d��/��4<���X%��#�Ȗm�����>���m��=�:\9�����s���(�Qp�8@S���nM��	��^�.͆��Ȗ@� ���ko�v��ݏNԇ����t8g�u�J�Ä�_����5�� SWT�p ېb�X@qզ��n�@�#�U�w0)�i^ĕ��w�WȿR"�C0d��X��n���)|��dO�$D���bMӽTʕ�t��*��;�*еO�^K��`�k@N	�G釳�3��e�����>�����}JD��S�b�{&*]8yA�9��A􌙉��;��M�c������S9[OY	�0�N$�R��zg�Rr�3���6�kX�mJ`3q�`%��A�O�T�}ֵQl~ĝ�F����u�y��EM�Ej����C1��ܼ��y�a�ܛ��\I�,�LE�}JɎ@ ޣG�0ʼ�5�������e`��Y����2�8n���9*Z��@P<�Wo���|�w>亶Ft����?����'��r�ZE�]@���-^�KFk�B%�xl\����F5f�=� �>��HP��-�D4�Ba1�#e�yK ��X1��'��o�Ŷ'Rd,�_�� ��ǭ}��gqF��$�]�;p��}��*3��\^� ��Ŋ�� �]_	��S����^�P.;w��>p]w�n���I���+��?��q�2>I�s��>_��٢�MWHp"�ښ�d�%�� k�^�<�ݛ *ŭ�WD.�������:�!��e��z�L��R1��騽o�O�Ța�����
$VN��Rb�(�\cC�\���iԂP�Cߝ���b~���6L��eY���>`͝�U
uZ������]�M�_O���}�c�"�?��2/�?�P�lb�%9g��$%"�i4fsMs��w������v��6Ք�/�l�v���t���?���J�����������߰��A"2 �ח̱���eh]�'?mgu˖6�F)S�e��-�R��"/�C}+.�ƴ�p j�ԋ�C��c��%��f��)ej���"�r'y��Ǘ������t7�����߫�!b��{x����߄<��%��<4��o?�?�n^�js*9�J^{w. ��e<EXq���*��3"�s�\�,�Q� �hE�=S��$g#��Sp���'MdHR�;|`�运$�`��H	��
�s˥���n��&i�X�m�������xQ�� ���f��Z��U���_�b�{���5��pfk<��nW3s���3X1�c�ό�I[�zu���EQ�������K���L+Z���`��1j
И(�z�Ctr$|7��>�s�7l�S4~EH�D2�0_���!4OjR�pX��e�EK�Q���v��k�$�yF\|�(d��p�n��"�+�D٭����ΙDs��&�2n�L=�/��U�[$��iS��ߟ9�&j#���Z�E�oJR�j\i���JgY�$�q���0
imHb{�z������gyP��%�Y0��<lq�fyG~�N>��"��`2i8��=8�uI���,�lK���'����R��[4��U��<K��Ы���7�nsW��+5�3�T���Y��r>߸��v����K����QEx��r��#���H�!0�*�f�h�d]�>���C�R\n��&+uJ�ǰ�PW����������N�9RL�\6A͓QE�#{�S�������o��jAt�s@\4��T}g�X�h��[�����fm:�p+<u�Lu�o�fŁ
�r�c@Y���\�:����tlX��%Jј�%:b��l�ܷm��x�7�V\���qܶ�C����Π�ӣ^�sb��&&���Id0o�4Tm�B?��n�I ���U-}y+:�s���F� ����)�S[�������1�c7Q�[r��lD�)��gȮd��A������*UhF�3�́��!�&}�t�� }��O�OAu��=��e���UD�r��ּ((�p��;ǉ<B�����g�Ta����U
�+p���h��^|C���8�/A��-���s5Ł�tOl���(���>���fB����lUM[�ͽ�4|c ���	i�Q��H�M~�5��A�NÐ��މڔ`Q��E?���<1+��I�6j���}^��h��? �'xD�4�{���H�R�^�@M�4�V~T�����ZI<<��Q?�xѐn�3�5��~c�����e���"�tK�,�+��f���h�to��_�\ [��ac�9��Z�s�6V��le��������#+�nk���|�� �X �U�
ab�j�~�I��MMu���s^;-y��u.��QA{��_L����m՜鮥X%-U��,�"f7�q\Wz���5�����U>�3�@���(�����P�z�-��g@�L!����$v �6�QX�	K�[[����>�C/w쭃T?��,�l��x�_������@]tp@ƫW!�6��g�p�ODҜN�e���O������nQ>��$QԼ8���uz�D����υ�w}"�.�sNl��]|�`<Ȍ^q�!ݵCÀ��
s �MU4yS�<�����^\�6������)ed��=3���r�x"�ѓK
������f�r��c�,��y	5�*��()�

��w��4 9%���@0~�Ƭ����x�-^h��K�}8әݼD��p����AJ�;J�Q��@_<��o�� ��uX���)?�D�K�B���M��F���<G�"����?�>�R�A��,p����O;�sV_�z��w���P���@4�L|)asSw�'�E3�UCXY�j���^rM���u�V��;7�����m\?�	����e�z�vߜC$f�?]6^=�&�71���w��MU*�%S=g�l��"�ZqA��3���l�"oP�7Y�v�U�=d3��V /ޠu���YӇ^��z����m�-'l���N/u����r��Y�
p�F��ߜ�s0�~RTՌ�l8_m~ M���X I�W������[~2���q��l��RW@�ۨQ�@��C��P�B+b�oݷS��Z�v<�f'��3
���9�n��Z�s�f\�ʴ��>Ԇ_��t���O���N�^�{�{ᔊ�5NS]�?I0��4�V�Z��Q-{r˅N\X�ZS�)�բS�I��w��$�3ow��~̖���W��ʘA���da��Z3L���r�2�j��u��]�)#��hC�dN7�QTJ����v��s�6$lM� ��	J(ʸIih���S��H���:k�^'g1�`��255~;�C�0��S��J�|���2ｃf� �Q:�����`�nM,���?�ё1^�A��"4��DƇvO�T�W�`�����\�1����9��c^�v-�*A0>FL=�_M��D)"m�8��17U=p<����c3m���T�����|�e�,�d�[$�N	�$����.��ZY�Mv�5B+5I�n��/{���EH[�gק��P�}ͨzm������ʹ\�����U�bp=2�} {��-ׄ(<B��0��9����1DK����睟w�����b\~�̩��$�� �����w�,��}�M��[��j��^*�^nH2��9��|�qP@��W�I4a��;�*CYh^W4�yV�� �c_N-g�@%[g�?���K���Lf#t$�iJN��X�y��B�<WopQ�d%Y��56П�}�%h.n��U��X�`tI�:���{y��~9�0*V���<;�]1Ͼ�Y���&���E�Ao�i{'��	��#����h�6c� �.��!�@@Ӊt�#�=�=}m�[��l,�[Y�a�u��ei��+��f�au{�e�:���:����Zq�����
*V��{�jՅ5��%p�U�p+�6�8LU���i"ͨM��S^�fvs�&3K<F�W�sڬ+��D+�n*�N�x)����qMA� #�X�~A\HmJI���'Dt�����2���p��~�#}ڊ?"�5̰���r�1�z��I��k��>������B�0������G`�]19�1o{KEJ�A���4�'V��wT+7��Cd�����[�`3�-ԣ�s�e�T俢��:(-�T6��~LT��C�s��m�Z8��ɏN�f�F|:G�Vt��R���q���*�]g q��I%������������|���ďKB*L�п�b�p��5[�oL2�v�jJT3���5�j���ׂ���H�V������_d��s�;���Tj��2��{|;��1��Di-����v����0�ϻ�%�Xǯ~���K�PUr�����yQb����0�? ��_Z���p�a=�Cg��W��㧧f�����f��/���eʇ%.P��r�I��s�8�����4�1��Â�Z���5|&��&{<9���'�g�;�k�q<�9��,9���SD�l�Uv�̬hv�*�D�v.Rkcy��C��q�)40tk	��x�2y���5����VY��u�m���!�~g�̎�t���bG���%������zZ�P�S�(��̢\��9Ҽ� ��U,P57� ll����/{L��q"�yd��־���J,lj%e�����tuNv�k�w�G_�k��fCA�>pp����CLs`������qRբ6_C�~>�8�8��<�9мH�uZ����bf�!�0��߆�uN��%��N᎐s5:B��(�AY�����cd�cS���yi�hv�g�yC�Yt�E[N/qP{�k	�a�0dv��D땦"9k��+��T0�Npy�P�j��T�~>����
V$s������t��x"�N�mfN��(��k��jV�	`��<�OL�ej���>2�����"��$�l�LO�EK2G0��癱�*�z��s�i�7>P������桼lQ���,�w��\���}~4�Y��9�| -2R���B��]�FX2@�v���>s�k@Vj2�?}��	(Գ[�NN�MS�5vK��k��~���޻ۋ�����	��(.�±j�U�*�{��]	졫��8��#W|�)M�)�p�k�A^�����2#���lm0����
{�,�,������\�2�]��KkЩ�ZBY����iDAÚ�0���o����L[�+i�b��{՗q�|�n��GZ���d �o`����kZb&1�f�Ǎgb��\iO͸��`�^S�چ��[�q9&�<���*�98{2�O�\nr���������ZlA���E�D)����Z���J'I�cp���Y�{��.ҖbǣvZ�K�Y��P9���Rަ+9��rMAL_��l�o���M�_�PF^��Zx��7NB�,j)3n6��U���K��c�$�=��g��*͎��P4�U.Ȃ>�O����W�>����_�����Jo{t���I����=��7P$k�{�%�\���p
KQdy�o[����]{��B�n{�@t�ܞ>�6�O�W�;���zZ&��_ш��j���-'$*y��0���A�􇜾{�n�Aj.d��(��4 H]����MeJU���SD�݈�瓁���@�X �Tj���i��4^Z�-�� E�HJp�ÄA�btW�P�i	�#�أ����e(�oQ���\��_�	D��7�3-y�s��
ɱ!�Յ��$�ƽ�d�/���7
Vt��g�~��s���q.�D$��B��]_�d8D��G��QS&�!�h��P�ov$*�&����;���,�-�|r��Wё���/܇\� f.&���	�g���$���c2����9W����Y�񫜚`�@��َ���m��Yd���O��҇&Rק��!�wcsD.K
��y"���;V�<�b�����Nf��s,/9��$N�;$��~sd�$+]���;7�4J�.���E�*�^<ݛڄ?�*!a
)Z�<-B|i��!�m�j�Q ��bsfDw���o�v�*W��U��ml�z���ta�@�rF*��D����0JlW8�n�Ǐ�o��3~s ��/h���σ�@�5��\h��Y6�lzތ������ )괡^{� �M�t	\�L�U�w�����y��r�=o�4t�w�d�-����\��t/p��� ��u*�R��~v����He���s��o�]�&��������U�Z��`O�K�k^�5��p�n-�^�p�B>{_�ݾ)��k��`��BU�U�$�3�$*�"" ò�!V�*��qzZi1�R�<?Q���JD{�`���ڱV%�;�G�)Q�nď�"
FVJѠ�+-�zCV � �� X���f��Cr�dՋ��rnu�T¹���X���e��g3�Ҧ��������!u�9w��A0���Q��f���=���V��C�����{���s���Cҗ��f��ܳ�5O�����e�Nf���}�
����"B�B�� '���(q����� X�t�I��y��~�y9�7�0�op��݂��,2�3�����(}M���7U�+&Ͻ��B��4�R��w��O,Mi<���6o�C��>�IP��mj����Uq#���S�i��v>�c���%��� ĘWS�时�2�In���w>P�id� ��ϊ����ic6���ʺ�As�pV@�K7�)��We�3M9�F%k̓؅��p�.���%4�%ʀ�����a�S�S����%Ȉ^f��ob�Ԓ������Ƙ^�&������;�o��Ԁ�݀�����W�fzA���ϲW�@A��������	M�&������Z�8}΍��zdƁ����B��k+�_C��CQ� �l{���8ݐ[�-�u}p~�тr~��n�!����N�j
zaH�r����y��
�����(B�n;�!��@A���K�`�wom��z����6#lD�A�k��`�8s�l 4���"�j��Ɏ�AW��g�;����:t�Eמ��7[��Ԫ��Mɞ�(X���Z�@:r�ӊ�z'�� 1Z�J��۽�a�"Ĵ�W���b�NpxF��f�awŠ�Tֆ�
��a%���y�ޏ5/�����bܵ��ʃ���	Q*�M!$J,5V�=]���?-V� �����h�ʤ���+�e����R���}؊^��$ Yg$��r2s�Zq� +��R0G�)���-���~�nY�s� �m~s$Ķt f���J	,�|?�zHz��3v;�J7�ּ�~J��4L��r˩��=�a�@�VN+��j5��r�3���p/��U����!�'�p��R�I�$�gy_�ټa'x<5�tp�7<sJߔV�=��`Y-+�� ޕf=;e��7�k�H����`>#�->��"���FUl��Á�q���.��ae	�Ե@ R��sb�l��?F�U��!��s��`�@��)�,�O*��e�� �hFA�)�����c٦�I�8j�4ֵ��lG�6ڵO��� �1�x6��ߢI�ڿ.����|ߊ~��+�X��D˝<���趗���7�5;�-{yF[@]��A�����{��u�U��L�m�S+�
��3q!% �x ��L���V�H?f\+��U D����TI���e��~����ނ��	3�q�����zZ�R\yN� �6�����沓5��`CL�~���d��Ya#�p�A�a��a}������2�I87��p��#�����d��W��Cz�����R���.���8})�r����Aq�nH|k]�{��Bj�������εK:z�+]������b{U_j�/�H�O�Xa����_
Ų�'<��Բ��u=,3&F�m>6�Uo2���FT�dCO�r����a���K���?�èDt{ܖ�k��L�-<y!C�.�<��e�-�]�:�.��[J�Y���}��Tð�7aT_�P'${� RxM�O~�$����5�4°��e��9���o�LxS�b����5��7���*C�L��»��:%"QҦ*'��e� )������L|~�n������L��aJ���:�X�|r�@T�'�8"�����>��jx��G��)$�<��#]�y{��t#h��kЄ����������#R��(&
��5���o�x��:�23m�D~�^� <��J�4k�-��B�������cr ����(R�U�@�a��YUᙸ8�']}ߨ �k���WR�i�ѫ���&����6�7k�Zr�aW����N�Vy8ѷ�Oﲅ�k=�><���_E3V����6���
q�ZtO����kt���6�����CǗ���	�K�s���*,�b���E���Ӌ���8���=�eՎ�An�ݍ��P #w�vE����_�MS��Ä?~��]�44����&��F
�7�Qa�>o�-p�$��v"��{4!H�Q��V��<TFm��úuDjp	&|P�]'c��!\�'@�3:�����v���}���X5ݔ��W�WY�hhm)�r��t��/5�X���S�7�P�Ǜ����n� oV�*�b�HDZ=H���%Qm�&�ܽds!�88��B���g�M����˴��|]itï�m����vq�� �x�'��g�c�Z���X��q����v0��5�6����l�v���Ym<�B���J�;W����J;<��v�Z�]��޷l�!6�8t՛׺�|�IzFhz��C����(���u�B��g^#��>8�^!��)7{E`��Y�����I�^Ӥ�5).r�	o�����l�H�e�kV�sb���L��mu���y�@��>o!�۸ꏟoS��Yh*�NB<�M�| �ǌ�s`���:%tG��g�f��Lbn�Sn)�a'�H���fD`�M�� "���t����ꗵ��VL+t��洓�_��9U�"	M��Q�LMw�y.�0P���Eɇت�	��}���g�*2�[L���A�3v���#T*�����I�а�� 'ZJk�%�6��~��m��E},kIL`\鬓�c������Q�Z� �#+�iz�b�QY�R���3���t���8OZR�=�E�����ú�h/�C�2���<�x˱�2�o�C��'(�Ew앲�B�@�-|��V�5�˳��5t�e��eb�t���x��5$*;Nи4E���Z����P4}����ZTfvG���u�2�w�S��O׻OqXj`�%x���L��<��H^ X�T�x��+��%2趵]�(�߂ ��y�s�s�OR�%^�ۉt�&;)�%�KQw|��=q���U�"�z�=�gJ:�����9`���:��RY嗲��LZ6�(��L�/�W�J.�;}�x�):�[z~��JK�Y����9�l�*̂h����:F�Zɰ��;zk@e�_��U��B�� DY�[ƀ{���t7f/�&T��?���Z��d�֦J��$*U��W��������2�-�Ps��#�4�
�8�w[�xҟs�A��o�Aj���O�<�ٚfv&��獬	V���{ѳ�(��rrn$�]�aWv]�T�S	1�%����Rh#f��˷oζBFp�ޤ��tm�P7��o��3�W��k��o�"BF(�d��Ĕ����Z��B<^_,HLN��O�k&(�Wd0�y��l��-(Yn}%G����-$�7>�����eT~�,�t|:�p'���&��h�ҧk����k���B��K�J����/z&o'2!ѱX
�>*�MT���J#T"��Ī2�\�]��m���}�����J���r����9(x'aU�x�Z
{�%��?`a�b�U��m�㟝~�PB�uj�b�$g��jj���B��L�{p�ｚ�<�W�π��x���^������j�������M�g��<��Z��2���46�r�X�!�ny&��h��RX�Q��RV�t��I>���~�U�ØAS�#�L�|��ň��/��B�B��%"E��ё|��=��ld'��"�:�Xr^ަ��#	��|#�fUʜ�|�A�$��0�(��Ĺ�������e�kq�ٺeԷw��T���UV^�Ҥ�P7����'��S�h �4��CA]ۺ :�ih^�J�Ĉ�x�[����l���l��DБW�h���}�[y�L;B|�݆�υpQ��k�<$9�)�:G�O��C��� r�F��%�y?$��Y���E� ��ψY�힧���W�`�y���e�9�-`�lq'$x�;hl<�0�t����Ջ����TW"wF��޲�ߏ3���58��P���*�D���,�[�Y�/�j��C�޲�׺�R��E�>�	��tQ�����4ZtSW��Q�1b�a���3�8���n=g�b۰ȇX�����ì�͂ b �bR�<��9c�9�ap�e���u�VE����{�U#R��G�����mP��AQ3E<��O!�:�;#D���p'���m�!�d�^SU�tI���aI���H4��[����1bo�j�|e��L��AB���b�ͽk6wo�2O2��N%9�uJr8>)���	
ީ����q�s|a�u��$�\��-���˿�K��8���}W_�����B2���/q��KU�"/<���W&�����OZ��H���T�J�ѱ^K��,1�it�ݏ�7z�̮=�21�c�f5 �3fz"��KE��/;r7w]���|O��.�A-ϊ���fU!���!p�#��V�Ĝ�1)r���j�#����˰$I�V��%��t���0�x&	e��R��e2���$�����{��[�z ?Rp쵄6�t4���7+>��vcB���>3��5����ф+���-B���� 7����DS�7�W�͝~�"��Y�KÉO���$}/��" ;b�fjA�1����	1�e��ln=GD�wq	>��������%���D%�dg�c��d���cF�j^S�H��A�v�;Ӯ����#��7��S�G���_>Cg�-0��G�+�)2]����~��h��6��G�P�� F�L��z���A/q�c�I��3�MEu�~�pӶ4y�!������G�8��#�P��[=B\�GL��*�ZF$f�MHo���tˎ��z�:� ��\�<I�#��C|��MQ�T� .qCƧT�Y]؏�(@���ή��н7�Wp~��ʽ֭��Iη�5��[.���K�@�E=V2�4�_��N�#�+�`7��=��9"@�uG��@E�CJ���z(�&���'�p7�K A�b����e/X$�-Cw*�˭M2�Y�b��2բ�,�a��������^i�Y�п��q��흏T,>"-�<�A}��to�q+�g�b}i�%��y��B=���&�]�=D�xs�a�8 xH��&�"��,��N��e���3��ϕeN� Gv�{i���
�1��6\�M�/��ݱ`H][�@JpQz���z�t
ns�ɹ5Y����0��.���e��E�A�����_�Bʺv@˫{�	_"P�ĩ=1�"����itŅ�lm�/�sfRN0y�I�6#rkUV���ާ����G��N6(a�Z��D��Ⱃŏ�wͿ:��s$�+{(�����>�!�����q*�A��=���	/��$�ڢ�Vi����&?�,O�w%����f�,:oiC>�˂�+>_��h� UK�8�P�[��9:�z�v<iD��N`���k}F8� [�~.�J�j�C�9���-{��g%]wU*{A��ᖎ�Z1��p,_��Tݘl˧M`A��縺E\��ROO���$Wa�s��@�*&�a1�W/sQ�l�X*��7T��me�7ido�([?w��EVaa$��I����m0G����Ԣ�<	ʖ�����b6��l�@Z��Kt�j\��;bz
������`* RHdae�9�F�����P�'�����p M��q�#	WHY� i_
�6��dФ�=s)Q&�V��^?y<zx��D%p�����`(�5-����S#����	ϭ��kH0�O�X���D��P�Q��4@9`-m ic�*�E����iq�)@h�.��4衅���0H�2ų�8���] W��=9��e�Yη����B�s��1�9�ole�rqן�XU�뉸�K�Ҋ2sc�K��?/���.���������w�X�pg��yR��D��=@r�IKy0��g �NB��L@9��W�4j�Й����t�0	!1���&1��~�
5�`t�sbՌ���.������6y��	�	��w�~��s�q��9+:M�(���K���w�[}1hG�zL��9H���a�����%���fG���j|�o���:|��R��σ�ᗗ3�j�QoV����a7!o��,�eX� ��W��z��y�0.^]��e�ʈ�S���[Z��=��')�U-.�?��/c;L��%�n�r��e,���+����G<gLD��Rr�D�4�.���vQ���y��&�4Q���e
���#YEo�R�Z O�?�\�_b�n�H�f�+��+&�� �DsH��@�qU�y��V��M-]GZ?��"),�#�sI���kp
�^I7�uO���ϖP} vo��3����~�\�1U�\�{��O��d�6�O���"��
����eИ�r��<e��J�0P~��MṚ���@	��$@��6���Ճ�|m�Ɵ&����1�0�	� p�n�5*[c�n������5+b7x~.�|�W��~�;eN"i��s8�h�`C�Q��;���6I��"9u@]@@'B� ���Ҙ:�Ԕ}遺帖�[M�,.��x<�IQ
 �AHj=�Ga������Z8�(�C@�K;|�D�J���#�R\����d��Y��q�!?Gf��V�����`.@e�CjW�_"b�1��ҳ�5��3�����{��L���A1q:1��+���(׼��ƣx�y[�a��Nf�":Ye �@�dǰu
 ��l]��zL�ť;g���g��g�2u@�UW'gKP��f!��ʳ��C<�U֞!�\��)�I���ee�y̎�j���bN�N�a���r͵�Xk�X�#�~r���M��꩛ﶘg�&
6.S�X�Z���[��b��:vz*<��̷�L�T<��VY2y2d���Y��K(����GP���X��
��eS3=~��	\/wNy*�]��￙�8�/���h"�qo+[���+QN��qμEY�Fsu��gE4���\�R �1Y��[J3�P����H�'�х����*��u,�^$���q�:�r#&�B�p�eJ=�7�*4�8�jr"�ߪ�=�O���������)�' ��P�S�a� �G:Z���:PG؄Z��ܹ�>#�,.��}���zb�]���έ+6�ߙq��~fX0CN{��7wM�=npE�;�Hˮ�hzA����"�\�������C�!���y�ꊎ��ۭt�\6�7/i���^Ζ��,�>g�q��~�*���u!�b�s]
�:����sn�/W0-��{+8\W)�i�^O>��� �=�a���T?\\ǀ�Z��)�o��r·8th���Pw���^�	�h�]��א4�w?t8���]׏��##8���7�0�%*;�_��?&����e�l���j�,n�G2b�Ts�y֩�y�	�����P�-�
���n��o�b��!i�u�F�t\<�'	V!z>�A:�X�CԚ)qiO��&���\����1�k!�A�}����A=��`�����\O�rD��d,���iGSP×e;\Wnt���!�ǭ������}�
f��R�+u�w��c)��.�d}�t��M����k��eun���x�+b���{���kL&|��N�|�p@�����]�U&CTvM�?�!��ǆ�r3�#
o�Oh*�E�]}7|��q��!&���3�9��C�B,���E�`0l���?���g����(|���?{!���DN �����D��g��C�QJ� �ɤ�`�#D�_4�&'~�t� a�+R���+���@.�����|� g���~*��*�n�j�u�%^�,6��&-�@�Z�,��|Y[�Ք��gjF� ����ς��Sɂ�u��dN}�U����?����Ri�?+ՙ��o�A7��nI��ݳ��%O���fzR]彾���#����#a�>���s��F
�����ߗCpۖ���Bh�ڐ� K&A���N��s<�'��SƇ*r<�_ [���ݮ6\���P�V�F�W��|��bCj2�e�h^�dg�M�w�N���Ղ?��G#o�����^mI�8*��p���ۏo"�h/�Wk{���\��[.�i͘�2_��L� �Bۼê�B����W���h`�ܕh�� e�1NZt���Q��E�F�aS 9d�߸.��Z���4# ���k��@�f�tZOk�o %=5>�@�Ҍ�6yb3�JDRS�L�]��=.Q���C��D�0�	h���Z����;��|d�1x:����*��A����b/P ǟ%��,g���'q��ٞ�)(.gDgȦ�kp�n��#.����v�n^��=E��/b؅����M;N��O:���ФP�W}�z� �kpfNy��8�0DB^�F/]2n���&@X����B��< -�B�C��&���L���0\ͬ��XP�F36Y��ˮ�٬���t��5N����x�_��,�p����6p7�TO���"�ޔ��v��V��*��m�jr@0�Bһ�0�ƛ۟��y���!��I����~�;φ� ��t�$ ]j*�D�P�����*k��\�x~�����p\��9m��J4���8zY)pu�R��U�CW�W<|+���u	P��s�wW?m�zj�ޭr[�K�>��S%��'Q���6��P��Ȁ!˦�H����0�7]�o@6�j!D ���),M�
�ytN?���s�����E���so�;����LkjZ��ՌT�_p<Ǽ��)�§�y�#(���R���;n/�wf$�O+e�7BN����Y���~�0
�.�hApa[݄�0�������9m���Q�$�����e����*�K��/����
\ɪ��M���VYe�n������Gg���x��3��&~�f���:U�[V�8z?���Tp�C��]W{��V4�[�
A�c�8�;N�����N�W��d��)h:�j�w�srj����;�>���
1�t�oj9<����t�֜$��Z��J�ɳ%�D<!8���ڤ��h���jv����4�L�ͦ���C�Eq����.{���z������\ޖ���k2������@�P|�PJ\v}��j��D<���o�l+E$s��i��z�^@_t����hΜAהv��Y@ߕ,�Q��w�&��r�:g���i���)���}.�����_ο��"��dͦ�5u��|�H]��{#�X#��\��Sl\���^ׇ�}�	���p^ ̓#wL���]c�	TF��=a��b��11ڛ8=����������*��Z�
:s�E1��
iv5�As%�87qY7�I�R4�������������v�qtPv�,����|�U���@a4ӝ,=M��,�~��/,1ƕy��;¼V��u	w.w�va���>O���w� ���s��D����W�/��_Cu�)��H�%��U��>�5FW+�o}�ָ�A��)>#��9`��8�����@�}Q����X3�NX��� )Ag�:�đ�WD���zoa�0U���&��ǜ���#��Jۄa���� �7֜U}�ѭ1�=�k)��L�9�����<(� ���+��N��җ��$[V��Υ�Czv�>��5�|�R��i����������(��sl��[Բ��eK�e(����@�bwQd7��ӕw�(b�H���CCl���{B'MD(Gމ��0Պ�Gvr��}2*b0�!1 ����Q���(f�~����倥q��럛^��҈3��NWyh����<�!��ݑ9�B[�z�\C��v��3����{�H�z5�dF9u�殁O�n9IB'\����׾�z�t�@��1����G��~
@�G*���YRr9���\<���#S������f��N���ӥ.m;I�	'�YԠ����2�{@���������[~YXR�M�lb�QXΐ7>���_n�]�h|a&��׽�/�I���~ٱ8J�t���}���L�9<�W��a9��yXa�s�ċ,�b�r��}�{�
��������R��a�u��X(���?�c�J�Z:4���}L�T�?+Nn4=^�-c{
���y�9�H�C
�c��a{M.�8��/6�1^۳e����Yn�Νd+�2�ì�a����HFX*O�w�ݨ�+w���a)�0��60&
q�b���Ï�Q�`���li_
w�:�����<i��D��7�z�.�<
a�.p�E��wh���!���	�0�}4�&QzfW�~	�`�c2�+���zu*9=�Q�u �{���)
��s2��/�5�XZ��QF�۩�:_f�!��~�O��G�������a��Yv8̧�����@s�M��*׏#��
�x���%��HC�Q�)G�a&hJ-)ҥ�L`�1����Ȱ��)�*C�W�u������%:ż>��Y�?��@�]^�,Ӑ�]�5BR�偳�XQ�+t��܄P��?���wܞ��bQ��h]p<]�L��Af\>��lH�xt15{)����$1�?�	�� n�A%�j���7�~�e���l��0Ol��p!T��O?�5�u�C�IG�C88���A��Ӓc������Z�~�qW��ç�5ޜ�4����4�hm1/]�G�� 0x0`gb�`�7��9}w�=��LXD؎p��(c^�^�W���8:I)}���Xs/��-�5�VPR'��Ds��@��N��k�e�7ڬ��>*)vu� !RC����[�w�c�\c�j���^!z�)�ͥ��[�G�{��jA�� �ĐҬ��9���2�Pz!��T;sw�<��X�;c�Li�I
�
��EE������=��Urɦo��$mC��=���_�[�j�#��䒅�#�)ܥ���e��&���	%��sf4�h- >L�»z�/ڧ�d�q���C�F~N�%��eVKQF�\����|�j���aKFA��*�d�O3~x+Q����2i��dd&K�k�yt���&�%�@!���4���������C��6]����r����J�!��Ao��S/I⣠$6k7�U��;�X��K���I�w�DjN!�i�-p�'�Wa��]�����r�7!ޓќ�F� �L;"����E�7����<�y^M��u��=�?*�yN��#� e�r�����HQ��v� ��p��
ZM����ʡ��i&��o̦�֯�WKυ��%�֯�6E��*3p@Ϊ���*��ƽ�j[NU�P"׋�$�ƽ���f6����z"2�6�&2�!Ot��L��g��"@�J��Ɔ1�_f�")?R�Dr�bLa\�aGJ��[��L�"91B�#_���C�XgH�#l�ʧl2G7�Y)d�ڥ6�����LP��?*��_���/��]�Ӻ�)���0q�Y��SDC���%�W((>[Q��2��`���8322�5���+��ҋ�7�u鮘�A5�V�e	��2���z��m�8�?cDd�6
S��R\N�-�c�ђ�n�����+�vΣ1�N�W�ٮ����LЁo3�Σ*h�ܷ�C��s|�8^��_�sZ�U29�ơZ�vyy�S�U���V���xO�_�5-��s�#e��h�-ؕ��E�8��f\V;}��V��:-�?�V�k�)b	vm�j^@��0c�Q�Ai�Z։�ݧ>��� ϑ��Î7x�z8J���78�T�� �k#�*��
��`���%�ɤ� �X�{=	�#<��^�	�2s�i� r�0�89sdV�j�`���]:�H�\7�$]��]��lM8\xg�$l0n.U��	co!Jn�y/��ᅎ��F�����l�\h.%r薠�Ӄ68��;�c.�{lz	Rg�����%9�fz��"���B�G�Co���&!!�L0�7�ʃ��.*�q��9�7F�`2#Z�8%D	����B$�?Ī�Iw���q~#�������eX��:�3��֟XU��|�~G�2�%���ə�y����7.�>��@F ���S����+H%F��v��ѩ�>���Pt�U,%Ikɞ�(i	7T�� ��Q�#q	�ش���[�M��\�����#P�Im
�b�ȥ+���z����Ljw�^�"H�W�2iAN�KWz����#}����jÃ >�gZdi��o�s>���R�noh7Q�d��\�#�t��^�&���}aSԙo����6wZWo4�c���9z��qd����AV<G1����ȶ�F �IF;N$	 v�f����Y1Osu;4��_�N�HFCz����>�M&��%��5�B`�5����=��ro����;�4F+��礊�<��A��]T�nD4@һ�(0���<��#K��	��\��#i��g-�E��R��u�[�1r(���("�aF�-���۾��+}��]n��^�_���U({aq��Q�X�"�%�tXK��x���8�?#`��z�b�F+tq��1\ےc�݅�N��!,��b�+n��b��]Mn~th�eר0�[y�,����*�-]s�����_p>,���ҥÄ��J}3�Nhο��QI3�M���ʔ�H>�@��L�<�'�L��L���0`������Ҏݐ���"����#��`ܶ/� d�mчQ
v,*]��\T��+u����/����;�k�5�}�4�R`��8����'���D1��p�s��|�:����o��e�?=ˣ�q��uuĀ�q��@���H;�Z��'�3$�|�I�������j����xJ^�:�B\.3�wy	�<����Oz�a)I����+ó�q��Z0x��㹂�x,Gǂ�K_��K{t`��<��:>���H������#$SL���&ioA/R��σ� �u#�j!Q10ܡz-��q�mβ����P�,j���wi���bFn�`D��F�V���?��w8J�,̫�>1����D�;�ݥ#U��}V�Oh�d�9 r�ߵ�����b��0RF�LUBX�V���/{�eGq|0}�_t��_~1�mi�4^M6������t��y�ฬ ����������Mx��y�̪H��΍~�&�}��q�Ze�3H�#�?n�UQk� �_ ���w�<SBͲ �e��z�稰������m�_[9=�W��V���P����N80�Ƀ�E)F7��'��6�Bpm�I��	���BZD���V�5�W�D2!����Ruz4u
B����}@�l��c�%�5 JE .�e��̓
ھ�檜�2au�_|1M壙D�T�F���po���%��`��O&���Q-��O�&Z�*��?�=�֯zvSzv_��V���&��&�?]��?��uq��>43rM�����2���5cr�=I�^��l���
��xeD)�5v׳P�*y�i�b�C���L�5������W�@G�̌X�]�{m�@�!�?��;�މ���+<q�(�[s�$N��|ɾR������c�I����U�~{��Ã;�X�tYE`�?.^:��o��,D�>R��t�� ��}w읃�Ɲw?�����61��v���è;IM������#�+�=�j ͹��:�{��@~�l��=uW��>�ki��W��-��,��x���4n����8$ؙi���=O�w� p�	����	�����Y��#�� ��tbF�ґQ8յ�)��Bf�y���LV51�*�w�`6�?���|A�/t7�u� fVy��J{�;
`g�����`eI��������������\;�6F�)G`˯�n�s��-|�r��^�����d����n����Q�0�`ʑewQ��!��N=���̩��3~+y��,���h��i㈊�������˷���	���m�p7vTKt�DI�˕�s�I� T<�i�q��a.4�P�|.tm8�W���^f{y�s�rQ���4y���0�D1#,c>�:�C^� ��;�
<X<:��4pu!o�P\i�P��W�����&v7�p�s� �O�gb�fJ������H������a�o#���b]�H��P(0�P��E��a�;�X7
��R�yd3�vIs��Q
��N�f����Eq�0���4�#Xس�`Fa����Ժ��/�-��'y�"�֕c�C'���*+WY�C��W�(C^��g $��d��J}�+�4�2�`�.h�2��T��p`���+IK
<�h�C�B��A�+�Ǖڒ�͆�Km]��S}��T�
r=B����U�4��d�[�V�=8��A^{�A��kc�b�#�쥫%�m�isI�-��1NT��s�p���RNj��oӗ���L����$�$8�l^��G��Aa_(�7r������QM,a�+����x�@�ȀWL��/����7cz��?����N @�m�9�ܱ�+�C�e�OC�$!lNMS�X��<����v�I�a`�W:����"5�J�!P���1�{�t���G��l<�2���5''d(T8�F��l��o��~=[���S����(�<*�'��r���Y�;�1���e�`�����6��%F�g���E�<(���k!8�7��׉����p!���x4&k��%�c���.(��lx/�5��Z�(U�B*]��ɀ,�k�U��w�?�{��b8kܕ!����� �↦���4EG�!��.��F���Xsv��V�%<�L����ݾb0ʚ��Y8��	���Dk�RR\�,u����J��ȋ|[L���L<g*	�;�UD�;�9g�f��Y�M��6�X��ZW�,����q��tQ�z�W��Ʌ ���r�E�ǐ��A٪�r=!"�%4����Io��H����A���3�PSA�&���֒\@¤�x� <Y��}[�cHmE�mŌ�ܢ�v�>P.����_'��[��h����W����u��X��l|�c�3@�������)}����W��i�S�j��(�ri� \�'�Pp���`�4*�p�~�,GS7D��C	q��7�O<^Y&��Ιt���$�ڴ��ngp�č^�A ��>9�a7��-��^��߹Ti�s�����O�	�#f+�� W�0�X��K�z7$=�m�`���£������r.�����R��b&35���`���z��L"0H|I��4���@���Dl��j�\al�X��<�|Rw���(S�K��7:�|m7~�wj��%��h�Tu��&��������!�͉U�F�g�,�̞�zvJ)��XT(���^���\7s$2�I�R@�xk�I2�7�7��[��ZT��h�A��zW�3�� ��ވ9�Q��۩��PS�|�ﳢ��O��ExA���@�ޢ����gJ;�>`�h(�TM�H���r��n����.ں�Z�.-�$�e���|7�#YYZ/���a�2M}�-%=�^��d���vV�}&�a������.ۉS]��<�`g��	��;��	z$%�4�?��`��֍�Ϻ��IObri�&k��[ES(yy���Ls��"[C,Ud��8�~;-����q�d�E���Ih�/L(�/�/��vL�w|�P]G�Δ�H���<��V���ǄE���ݸa�	�B�x8xg~�v�/ x9ML7������4�(�%?L~����X��y��0H�p<v����� $��?�y�ܻ��Rn�b�{z PRS�|}/���]���5��C��2!���$�>�)I6�ywtׄ��qc�^3{��=E ԜA�H�L|�j�W�%Pb*З�"���߿���E�~��EL����B��kT� bs�,��EAw�����(yZN�D�ݞ.�<F괶��9FDX�D��F(G��ZW�N�-��S=�.�4�PC y�Qq�h��J�,/�W��Ey��x;�,)��lB���Iq��o́�4��g�D��m%s��49��=���Y|�e`�o:�;��;�W0����(t'�2؊��K�!�/j~�k9�ԁ^gxI�ϡ)G���j�0�;6R�Zw��x�/�!�~/���;����V��gvP�|Oe��w�[�3�����e�p��� )�<Zl���N���Gx�혶=�<f�[;!f�	\��?3>٫n�qO�a$B�L�^��M��*��o��:��Zށū@?u�ήk�z���.�X*9�ú����Р셖���z�uL��7�ϚM�gꋦ�9�H��`���7�!E`O?O.Kq�`���:�!f_S�t�:>M0���	6i�����3!��3�@4�f&�m��WX?�j�jAʸ"���ix6X��6�}�{CP�A���r��w�,,eo�����ԮVݵ׫������Ö�y�!���H+A��I�q��%����=��Ľ�J�m�=��o5��z���r�¼������qk1Q��W�UmH�ӂ��p����mY�E��%��sZ
G�k��rz9��?�5�t��k�Ů���630~o3�c2oj�G3Q��ŭ�qǻЗ��e�1r
*=Z���"���65���*q׳Ca�z�cH ��Upm��GlI�@`}>�?��]�!����M��p�+k.TNNo1�G����[9�a_]��M�]^��0���N�_&�OҞ�x_��裞F~�D��U5�[�8w~�,����@�BY0e�+�j�\/?��w+��9y�F7���b^��-Mvٝ�&��/��aL�m$�\���
��5�]�G�[�p���s��_)�
�U�(GpY�ٽJ� ��,o����@�c� 6���A�Ʀ�H�Y>�X�wg,q���E�B +����We6}<�9�!��Y�f�= ��9�!n�/T	=�
!]){{�ܽM�Q�{��K�ұ��uQm�m���=�{��*�2QV!�7`���n����[ �}u�$wM�3�A꡺��
��m��u+��3����+��Q��B�jB��u����Q�=�GMp���}[�Mr�TK���àt?ކBgE>ܦ<1�R���߉�pGf�ߒs�$W��8	:���=j�����H� �M��[��s�G�1�� �XA����LĢ�������γQ����dCIߓ'���K�SJ�[%"�6u��?\����b��P|*X\ó����c��3����A��(���<"?���Z���'C�r����&8VfgQ��u6VhƹqR�����9_�D�&I져,���ೱ��z�����$�0��,� GH[H-��7�T/�'6fa�&�µA�O����2��M��4��}%� �(
$%���Y>A��:Ք�g�ubbv����|0�O83B���8j�T6��SC;0�pA���p9���^��6Y�Ą=:��F��ɞ��ck�$"s��i����K4�Аp�l"� ��)�x� ��DZ���W���@�Z!���C3=9��	J��:J�Q��b��[ʀ����&4q{�C���e����a#��h����ZKS�tz����t�^�����{,�v�L�#��_A�ISp�W�G��8y`��5 X�^
U�;�h�RI�6+} 0̹�GSy<�f׸PZ]��NEJ��ܯY+����j��${�SC(�B�\ks��ۓ�/U�c�dpC�g:}�}2�r�=��b|��-��k/j��e6�%� ��E� �������]��r����ut	�5����)uYS�K�[9�j��`>2�ɟ��c�yQ�������h���Gh��$�:���u^�s�1�半`���r�h)�*�PG'�q}z��p�31LTŭa��P�G�p���W2F���|�.	E�4���<���`Z�����i0'��h��X��e�s���q��G��S�Ӗ���Vbn{]5à�|SX1JF�A���YRC�9j���X;=��om�OTʃ��$����z��w�zE����FA�U{��!ѝ*&|�膵a���EE�9�c[D���
UJOlD��,�8���G`�K%����P��`�C>�퀤�u,�n2˂AYy�x�`��[b�����jTc(�k<�
����=+U'�vRW_��m�TRs����\�/u/�1�҄n2�c��Ӄ3��L�2Q�4o�K[�2>$�7ʕ�=����:܋J�E�'i��� �V�+$��h�`.�R�r��ΒUaA�֍��Ե�D�!{��4��ɪ�ꓶ[�������-���*	��Gb�[�e�y
$���̎c�@��t�.����nJ.�å�Vͮ�{H8q��x�չ���Ә�8�$Lyf��S�E�Q>.�>SyԞ|��Knv�[�X��VЂ] m�TH�g�y%5�6wQzi[Z/��-�R����]5��ҴDK��ݺ�j��2b��s��h�F�}�T؁&���S��(W���Vfd�r܄�#�l�(N�3�^V`��;6��2j,C��v�"���ٔ���c�&�������O&1p��>`�RbAro��~�����SB�����V);t�^�%RGv�^�滿^�i�⊟��1��N�ŝKv0�X�F�q����ibM@��^E�|����d��9�*�y7k1��AцzX��^^���P�b����m�����-'��J���O��%��H�sMg�[m٧���ԗ<I��I۝�2�`�T���ע�|�<S��s΄���+Zv�M�oD�~nr���dWx�ܗf]f�ʰ�rǖ̝�q�d|e��?�F�Dit���.)O's�@�;2"���o0�e���xy�W
;860/j��]�Ry�C����4�-(��\5 }v�T�H��� Z�cH!��R�Л �:����n�f�f��j%w��*��TCكS.��w�q؀����3�Z3�ϔ$���Y���1Ë��tĸw���<���@�@�1�{��XU�xhJ�x� F�s$�y��&V���>w�5�' �R�B��"����p3���;U#�x����oj�dѦ{��~g:_��{������J��O����fq}7-�)�7��Ԉ �S4��;�̎ v�_�t��J��W8J5��w��n�{�f���}ε�a��F�L�C��9ɤ3t�`k�U
-��3�`�-��HA��f����X��)��yO��9�o�l{�DYEɭf�۫��|�ˬ�>��4?�-E4w�z)[`���L�ɩ�8����F1%��d��܃k�ҹLrB�D�~�<K|� +Y�䀮���D���m-����'O0�#V��X��oq�ؤ�����]l�nJ�3�����m�JW;��
hE��b�Nٹ�G�gn�q�j���qY���>�����Ƕ��g@Z��.t!-�3'^�ṭ�3�{����ԞO -B뛽lS���>P}�A�i�ֲa��������_�>0�dN�iT4����l=��2�#����4M�ym����@\��$����(et ������C}�Jj�zkO���&O�5�k�M���6g�M�D)��!�bP&*��9�?�V�ص�/ڵ顜�9��y;8B@f^����*�F����ī��#nߝ*��i�nLwdʫyu���� xfd�T"���Q�4?�����H�(a�R{�{�d�� ��������b�[�Mr.���M�ǒz���Wj-X�pj����P�D�@��CK�r�3Y~�P�_��ڪ�m�lg��7��K4@>0y"�Z������n�P^k�}Œ���P;e 3��
=�E^&��zzv�[M�D)�f�pXHxX�T:�yj��v�U'����ej����ku]��ݣ7w3�~���n*3oNO[��R�z�J�0j������S|������tkG\��Y`�}�e�4��^�Nf/�p�Vޫ���+��S��&MCe� �ho� >2�~��ެeٹ��]��4�H�E��Mt�%���p��N�O�I<�p�H��R�"N�`+�Ј�29�"����`��tC	��n�59�:�����7x ��kA�FjbҘ���ݸ8�7��<4�ŜQ|��R�Rk��k���2l_RM��=PerS�Z��3ds:;���_bDY�YASo�eʦ:Y���� �:kh���8�>�����1��>��4��w���+9=�3�NA�'IS���=tJ�M����=�[�����[��;��h����NdE��a6�n4�y]��Xm�������H\���	�p�5b��w������7s
��րr�<���G�&���f�㗪ST�̵��T�_Wp��_�t�����w��1���)���5��쁪iϺ��4�e�J���� l��ڑ�����ؔ'>z�I62�fjOW�s\O�{�jS@auu'��!iD*9+�A�\��o�� �������6 ^�Ɋ�5���`
��l���Bώ5os�m�`��a��&Br�i̗�}�X��;!���vf&�xe*��~19)��'�.�
���{�":�Zƺ�d@j�&���8���{����%�r�´��;�bb�t(5������4���Vq}f��y��˘�RZ��%�ck�
��*�#�h ��: ���2(x�)���K�إ5&����m�e�L�gH�RX�.�p�yG�!fEۂ�O���uZ��kD�M�ؓ�x3q���RL��S�+�������΀:�;y(J�(��*�-H�T��&qr�v}����k�[7p��)g-H%����96s���C�4G1�����k��g�/`�b��������_v˘���0���3��xP�)
#1������c���`״�s�1�6���j�2&���
�"03�J$��H���8^��[�P�B�����J|�Xɦ<���T�P	5�O�ۣ0h�T���w�هh�|Ij<]Tà��y5���؉��C�r�Ƨ�#/����T?
y}1�[ç��9��3&iy-�G�yG�P� �S����eY���L\���O��?@g�\�#���rvi�7X�`�ԿB+�B
;�$X�x6�G�*�.}?��ʺ���n����檴ٓ�� ��D�2�7b��-�����m@�|�1� �(���6����W&�ի�&��4'����=/ȾG�
$�kŢ�ު
�>r�ʦ�A&�L���S��|S�[Å�l��k�jv檠�]�B_2Xą.��������?���1��rf���tAjyƱCEmc-B��7R�`4�C�s^G�:�Q(g/��wF��sz������3�6�I�wI�Q�)6u-7t��O��1�m��5�I$g��A������E�����C�ޘ�c�j���v��I�|�j4Vy6+>������t���6b��o,H�[^k�A��*�Ti� �j�e����Qt�ԝ���l<!�3�Q��\L���u5k�ܵ�R���[���O&�Y�?`>��%+܉L�vAe�JyOO]�&��ܼ��������bszX��E��H\���+�ȩ�����}�������ִ����$�{��$�$�tY?�ܬ���(R�Pu���"�뭕uwY\��w|��t���
����D�4p�:Z*M�6���ɻ)*dR��[xe�p��<&^jHU���)쳀D�d�#�{!�Q�F~wP��k��3���qm�P�f�G���T�����(���a8�@����3,ǶX��j�_����;�BR��rT��BZ;;��-��ӹ��9�#}���r���e��l��c[���DFu����RL9�H�|`W�>TՋH����0�"�S9ӿL�<U.w�-s(�U&��b�P�E��1��R�cc�*�EZ%2�&8�wU*� D��ވ���]�R��Ln�����'1aцK�(6d���d���YW�� 03�<��f�ܹv$ЗѢs�����r�A��J,W�`>��������rފ����'��i�p�|w�2\�Cw%�c�_L�=g<�`��"kN��)6u��d|� �:wI�
_ݑ��|�ݎ$Ɍ{�Äb.'&@K 4$���M$s?��P������$�q�����@�=`��5\���A0�������5"I����)"W��{�a����cȰ
0K]�v�w��t��*2:=a;�*}3))���́U�m�Lug�ll-0�������3b�E���z��6�@OK�?>���O�'�C�[#��r7>���B.䍋p�#�_ֽ�H�4'��,��:�Y�]�D~{-�Z�F����/�7��	�wU��$��=�D�����	�z��6T�h�V����|ddQ����c}����G���5��W������ǽ�����@��M�y�N�U&��jQėT��v��pd?|XrN_3�r�ZRJ�\�|g�u��Z��9��h��A*Zڬj�(!һ�;�%��T9o�ɕ�b��O!�Y�+���2�o���Om0�j�,�=Vx]1�� z�W�Y�ˑ_��\��Κ^͠�>N�qN�$�;.�^�bǾ{�����hՃ�!@P� '8h���EY�A�k
Hڍ)�I���"r��4�����O\������; k�,��6��;3M��`.�mә�cS᧨�=zJ֪�+D�垔��[�֍�)�|/eѢ4�d-1�@W�I�#}��7�9{=�B��[Q��m�Л�4��9�p�7�r���`��[���J�7�XrĚ����sC�z%V ��,�|<���x�
h��ӽ��;\yZ���}�-��u�O��L���r�0D�w�j*��I&��9DSG�zR����'��N,����hA�J��cr�'!j��3)�2���j��
c�ˇ?9��^�^���9S�@��ǡQa6��҅�����cA�յ�ߜ���>���3�3%����r�FY�������!�k��ja7�<��u3�R�Q3��~W�jO���>F���]�$zl�L!Ə*r��4��TT� ���k����լ'��n�����:��\�I������i�MV�lb{�q�,�Y��fQui���G��X�jU��6�խّž��r!S\h�&����]�"kX�9a|癴���-�E��Σ��c��¥��f�j��6�>�U���3�~=|�C a�KX�Á�`�xv��0������t��*J(w~�%�%v�de3��$y�7=:�2�K`|����2��B��F34QDv�=B!��!W�1���e���TF�9��n���h[}���4pM�/;@���:x���;	��q #=�~����|N��A��xx����?�<#�*�v��/Y��2�>r���؇w����]�s!�$]v�g�&E2Ej�1�Nu�6\�=2�j>�&��ߥiL�0	�����W�����k]B�o{9�⫻�~��֯�v3Cq�"F[�\�HPf�#j!����@�^�@f�k��D/d�T� ��<�K�[ޥ-�ؕ�����)���E��4τ�w�8xsk0� ��qe�m��N�՘twk�q�c�>3P	�ג��Q-,*��+X9�#�y!��xQ�J�-�L�7f�m�_`f�I��Pzr70m/cuXd���8��a�6�V�LS+�6y�'uo0-�K@@�8Zmx]q�9����*�z���6 �7v��8���O�ݞ�����~fau�$X��V��fn"J�8̽�'�E��b�5�歞OQ>�j�Ok3ۙn��,��� X%LpYPG���/^lo6�H�PHϱ��42��0�] ܪlǉ��\���>h+WL��wV���qdt2��a`�?]⎶�qX���a�����,�����a����O�E����I�-�:]�,U֬�!E���I7y�1�	g�S���U�M��r0�%�w|�׫%�C����L�=q��<]S,M7�[16a�2��zï]�g�nV���y���ϩ�.y[��q�L��Tg ?h6J�._3�6`:�I��zkl���h�A����'E1�4�Z�����L��wnǐ��[�j��G�������'�a9"�iV����G����G�����;�V9%�@C�������C�/h������@�F��uEI��8V�
�H$p׊�95��29�BD^2u����؇	ܞ��}^�9Eܡ� S����i`=� ����ڳ�����U�JWr��Yd;������-�ӁU�p���PAM[5G(������+��f�B�4/Uє8���8*����(��օ��6i�"�u��@x�On1ctA���19�4���^��@��5~0~��<Tt�5�1�ɓ�Ds��}h��r��7[͡�J|GKn1Ps���f����\�e��`�,x\|��Z���FD�"�r*2�k)�I�V���"�Ǉ@<�~{�FixR�>�[�U�|Xͥ ��(vp4p?��f�io	�x}��f��0�\gn�wR˂M�}\)
B��M\��S-4�T��b�]�0�i�$Ǎ�ۓ�0j!�EJ�q���vQ�ԉ>%R��`|��B���1V�aZ����'}("_Z��Z�f�Y�_�.�^j����e�W؎�D�|3����7�%/�����+M��	�Ӽ��B뱰C�t��WV����Rt�Е��"�����j5f�vQ�g��G���cq�ȭ,���%���
;���iў1����8צ c��c�"�O]�5�ḕp�wF9��yc�t;��~Fy?�ŊuY4,)3���⊾B�,2�y�������$��k���S�P:5cc�5�����佄�=B������8 |��܀ԛ�>��݌w]��$��|�����J޸X2��IնѳJ��S����V�4;S7�[����w���G{59�W�'��}�~��3џ�Am��D�����v��.ָ�l'FK�D��,���~�wf� `�N�f'y��3^�?���R�M�����k8X��B�5�И���ґ��69��GiQ�����5j�ij����Ů��A;@��X�����Nc��ŕ%��$d���j�'W�hI��ˬ]j�|�Q��MN���@v@�t�� Ͼ"je���Y��|����!�Ku]_j�꿃r�{*������� �~�zu�m$���M>WuE�z/�Y)�r���-f��"h���������[v�%�u%OVEn�)�R_�P��*"!#�R���8�I����7���o������9���'g�p$�eު[�M�3D�񇐈-"ǿ �t���bڪ�?n�����kv�x�,�Ř��� ���vo��b>h9|����N1|%{WN��Bƌ����nW�'�f^����^;����qX*rp'J���i#j��� ���1?�)��Ù+}$���Կr�DH�p�Q�f��p�Y� ԢMdv38-@f�������2W*A^��窅���x؅���c�4�����[�DF��:9O��[��6��.p��'m�0R�-�p&����h4*=��X(,� �G#��Ƈ�KO!�eQ��M0S�~*��ʯ�(�co�C�t!J��!�e�?P�T��{�#�����S��}��V�� @wd���UU��L��M��V�L�G�\���ؐ�Kx*�w;P�!�ґq3���m�O�d�Ap�8	[��d��͑S<�*{߻��>�P�Z`�"pВo��K�B�ˁ�~������N]�l����/Y���GmUd���`�X�P�д��\H���d"x:5O�m��S�Y!��m��Vm�;�Q|~���d1�J�+� ���N�u:�u_T���^$��I�`,/���{"��J=^9p,n9������h�;����\�ާ�{r$�Ί�V�r��aq:�y�-��\:�6���{�az�R4���>QGcG���*ۆ�9G���s'c1�DJ�v8e
��&c[��#���N��G^��Y�E�1^�7%&��,��ˊ���Θ�_�?s���fu�yguși��mR���	��<TO��ۧ�[�I��BN�6j�П���hW84�ܾ����uJ�t'KszQ���=cp@:�v4 ��82�HuaԪw�~^�_̍��7XB��nm �J9�A&�� ��n�k^����/�/!'i����n#J,�0����h����쾲�-��/[�;$R�{-X���粉l����<$V�g!`����#���ݻd$p���y�f�HbI� ñ���-��*��5�U+�E<��\�9���"Mu'U)�%�-L��� b�2
��@/G�y�$����y��1����s
K���Bj�F����?°�,�E�}Y��-�2F��D7w3�1�/H@��zě���v+��L�' ��5�qy�n��:���u`�NE�2�q)�#�5T&��&/�Q�V�y��NSjp��'��V;'&Q�
1���*5HR�S��u����;-�}�:�H\�hl����W�A�լC
sL�(\�*(�8^��vu �+
��bWUg�i�cP� �Д��{��w�9�Cq:�%�W�>c���߀w*�]ߌ�_B�
{�C�=Ad^V�cO��;���5���(M_[b/3 �� ;��T��	p��Z��,]���?9�KW�CIҵ	��;��|����}4�*�JUD3�Z{0���	��i�!V��zCΏ�}����Ʃ.�ϒ����GĎ�mi����j�U!�L��r�^M��A�c)\��Wt������<�x�Q�L8��.Y%L.���e�@L<�K�	6M��~n.Žא��0b�(��>'�����*�>_Ȕ�8�t�L+F��=��6x�gVW�"٪r�-��Nv�I�:`�4����z����ך��+^�E0�hՅJ;�r����JE�{,���8�sh�o$t��6Ә��ڸ��9�Ze�ʩX��,љ֚��0�Y�T����A��6��ތ< �~F�:�Pg��s��M/��l
RC2�0�Z� ��8�Z��P���hf��d���MQ���+���dͷ0�O�p�b!��8~9�ra,u���
��0_Z@ ����������~��L9"]ԙ$���EpX���9��L>��o�A�5�WFv�l5������|�I;^-Jd�!?"��z]��u�g��5q9��Z�[�b��Wͯ:�|���b��c��o���xys�/���P��I>r[����{z��M�x8y���2:�u�d�S��^Y����RLox�n	ߘ��5ckhG�|yzÏ}�g
��<ĉ6�0�s��/�BvT�UѶ�� =,[�qV�M���t:�f�j+J~{Ҩ����R�X�WxL����  �IޛK��,���&�<������ˢ�ՠ�U���}g�ŝ��0�v\�.6U�h��ķ��孁a�>�5#EL�2�Q�"��ކ#ֹ���=􌁥������,��Q���[4X�(��U%O.���F���A���r����y%��i;� w�>bөoz��:IQ�?���D:Q���!K�n�]ӓm��p� �	LTj�wg��(��M�u�GVo~�V{���-�-�eL,�	�s�5{K=�?�A��{ya麸��M5������;i�Һ~,>w�����(�����(��������1��ɛv�������Œ�4oW��������-�� B�l�)�z��@��q�)w��i��A��;��� ��J��PF�X���gu*6N��l��cKu��-�je�4�]'�ۤ`�N�9Zw`�ԟ�G;�e��YԤϿ���٩���o�%��-k_�BM����YA;�^�];���Jn;�qcT�c�<�:�#~��C��ʤ7��sB7:�+6S�Ғ�Bq�=|��G`�`�WUϸr� )/�7�S�l��l���zP�QZ�����z^���
�N�X@�&ԫ�ҳ��H�_>7�أ��qZ������W��ߚO8��̾�����8-Or���?y/��gA�Pe�^O.��4���s#GY�[����ƥ�<b�cĲ���uo�M��<^�!������=HX��e�C 'S�(<�_��|#&<
Ϋ��G/ Y�X���9S٣₏tE�JK׀L��Bp8`~�w�$���s�Z��~�}�"XJ< ��'c��@�c�?z����t��QϮП��������>J��N�:'�׆ɥfZ�����:�U9��qo�{��A<s
�w��:�@�����鑊	l���m�-XW����?{���sιe-I�<�z%�L���lO��eE�l�5a�dA�RWx�z,�Q�.�cm`�����!�
����=���
.ј˩Yf��Zw���ٯ�̆_��n��8�Xa)�_!��T �I�[\���#���<b��Z��}�.k�0.@�	�Ϫ�Ȩ���ε��Z6�=���gUٳ$*�~�Z̈ɏ�����lZs�������N%��1�d���(��_��uvw�������_V�&xg<�Ƹ9���L��������
��2���!5�\��9Z\��\ć��_R9.������Bt��%�EPRG��˦�P���G�Dt��Eqݞ��!�.Z�l�'��d�D�������[�ev�*"G��b��A�+Т
�#�\��z! _W��j	��(❘K^���ºl��uOL���>�Ԩ :{m��C�~0=�i�ھg[��"Poўɼ���{0#��䇢�Mʿ(R�D(Z�}}��y�+1_� ���8�� ��)#س���P�#��v]r���!f=xMxS{f�]�Xw�&�u��g�6AH|�y-��L���G���V)��s)Pm?�{�E�s�{f�?���f���	�U8t�5���,�f���Bwis<��?��cl�^���DȐ
�3t��ra*���E�>��t�4��4Sħ0d�lkUo&�ȇ`�}�d�C��	�A�h!���GD¿[|��/PN�.{[�C	h^����p��}�,�f��h�_O}o�V���iQX��s	|�?���>�\�7�*�׵,�s�6૝�yD*�L�|�jnM>����x^� ��b,bP�P3j�/"��9��?���}��S����l�E���`�f��~Z����02T��w�,%�9������Iᄳ�
,����%�dI�ݪ�J���Z1&/�-��83�	�X���~��|9�s˭�K.��k:aW� |+6��
���h�/Q���4K�m�Dq��w�d�'�W0��xy�����/����إ���(Lh�p={4f�������JH�"�ybp����a��Aq}V�(Iە\�:�02�ti�l4u�샃e��6�����E�M�����_�,��)Q��d������=�@Kya�Y��>,T�.<2�+@jV9ZUث�h;`�����fU��Eu�8���5�(��:�G?zĸ�	I�{���E����4Z_nY�^:?�a.�W݅�[��3Ã��(��/��I1���;R�P^|��j~�kK>��@�ᣩ���J��tl�t �* ���g�
��위�����?Z���gA��h�-�����FTZ`]��	j���3�H8�*��\���U�儱%���voMm��� 2��@���6]��_��Oq�8u��`*�&�������������Ә�S���IE��|]ٷl���� r��3cY��{�%��p.Q�z)9n[����5Q$��$%�f᭔jdi��<��!ƯuZ�~u�w��_�GEa{�-M�7w~�'���<�����ʈ�|X�w0��Nb�n��X�b����R��߄S�AY�]�<��*���5�׀�/�т@&M��>x�@��T��eŉڟ��,��2$��{8�qsQ�"��4k�tk�v����adE�j?�<�h+�� ��7��J�� }q4�*8?�]�E�H��=KĞ��)�O	��bQ� �Ș��$B>j��ϳҼK�Y�v3e���ǭi��&�q��N�������R�_�^��ʢ*-R�$̓��_�)���{��)�2�<�W�˿X/��6>nS����X�wo����|v^��[������0�+����*z	\��]�&��NRK�}Z�-t筕t'����h�w�zV'�F��3�X�9s�>�e��Y"� ��L
(i�{�i]�-qg�>�Ւ�E)��*�:g�-�G�u��>_@!�<�!f�|�'��9 K�Y���Aa/�#��)w{h��{�p��sS�a�cV
}�"_�X��&@0��H��=�$	z�E9&��ʊ�e?���T�_��g}b��V�dG�H�����w��(CT���p+���2u��+��G��� �'=qFٵ�.m�y�O������gS�-'hӥ��Ί9Lc|�`�� Z&_�nv�4]���=�5�
�_Wx�m�!D@Y�����_�����d��-�a$z���?�w��J�t�"���jM����LW�ξ��N|D&=9�Ѩ����]gZ�KQ=��
w[��\�ot�m�8�V.��2���#i6d����c gDƍ�p,'�y��� A}�3��M�1�6��GP��Lǐ�����W��bF5�Ql�l0m����h��a3�$5ZjpE&���j�"����\yY��}��R�F��ޖw��a~��:�ӊI����~�US�}��F����tD�6�wU�`�$���ύE�����&�F*0+i�&�vc�Z+%� �י_�v�Ջ̲2]���wP��k���$����Γ�±�*�|\0 ��EO�%�8���m�M��̲1v�ڢ�	��g-���Ȕ@���e�O�в��~Q+}v_�rwJ�R_����}�R+�����>���ഐB��N_ǧ#?S�Ш�:xN������56�@�4C�JG7�C�l���[V�٪�)S����-���r���֨�1� f��q�w��4������9�b$'[5T��+$���D�-��N?��)�%oKW��/���c8�tׄ����T�ەsL���U�gm.C��g�1vK*��m���z�K?F��zG� ��r�f�� Px�0eu�B IZ�$�H�]@� 4캫��F��R���L�o?����;��σ�Ƀ6�	��fk*��2ˁ�K��p�Cܔ3*wOq_�ka�,2�ÿ�NǬ�%��Ƽ)Z��Q��}֢:��M���qM�����֑2�jU�R�p��0*\X�į��3��ś�5��[a��7�`�<	�qcNEO�K�Y��m���E���2N�v��M.�	{1�L�;�P�Y�?&�4�?6�3p����Q��UVY�Q�t��8�@�`�+AK�<��&_"�����S��x��g�v���2Z��X(_Z���{[��p�&����%bhL!���|d=F>��[F�:�NU���D7?�����S�Y�)$�Un�����E��~t�������쵅���KH��%Y�����O��R��PP��Zc�n���"/Pę$�[��+d�'�ם]�/??C�[��Vqmx�|�]c�R{ę[��0i�~C=��=F'�����@oƑ�
�����8(N��̫_�#׶���A��N�3GD�.Z��8��v�]J&\�g���8X��.}�9FUFCL:V���o��6����٣\���d���Ž�N�W	�l�उ��E��2����T��L��3�.��_��-�Z#�dD��7��Q~s�}�A�E"�A,Sq}����;���h�i�T��^CX T�I?�U�sYăM7�ݗ��#Tb�CC�hh� Q_�M�.^����.��Kzp��1�K��dA�[D2��
�ڡ�7v�	��4R�]֝g3|���:K��7��E�C�-4p��+�Y���'A:?��`~��Y��s�n>�R�d?�`���{�xB�T�.�_]�Nۊ�HmU�]b}��d�]G�i�"�r�1�����{"��(�WN���W:�9�����E0}'t(Tm{�\p�)�jDa@fnh���T��U\Ҫ�U�����x�9T��릁8��r�����(r�MBч�mD��0��_�^��%W��b����4�Z���EH-Jvc'�]S�3���PR�WY���AiODC���	�]ar=*A)��V�����++^�

�g�un%*�Ң��ú�"&�Д�~/�AJ���-'����"�x�2q�s;ې�QG��m��Ik�q�h�*e�%ee�@|��w��H�j�_.��o�2���3��䔪����R��G����^|.L,���P���5�T��
�kػ�;��*�r���"�54���d�PCI�1�P��A���K;F�x�ZG��p�#F$ge��q���24���(\@�\�j����Jʧ:b�v=1��<t8y;�n�����<���������s"��vfڴ�0%�f�*�͍�={����H�_(z�����W2(%��P+T|@�������p��ɖ.<��S�BGHL��2����;�`S��p�<=]��DR�S�t���Z�j�@���D[��8+��ր���@���W�X|81������ =����5�ﰅt&�|{,��8�ҹ���ӥۮ��/���q,h(»��]���ްS��t��2�z<L!���h�Ø������(�oTo�f��$���ZR�ص�MD8����������~�y��c˴�H�;��
.V�nq�?tSa���+j���O���o�9��~s��ׂT�9E�ꧯP�������lY���}@��F̖k�N�tW�g4ڠ�P���%��:��Ǟ5 69����V�\!�C�h��]�H?K���(��T�AR����D��[;��nx{D��zn^R������L�����K�ƊGm�7g\ ͧ�D����'M�IF�/&��ᚆ��SV	��O����}#��H ����Ws!�A@	���,H73��0��������8b%�;��.�Ί���)��i���7xU��ϭA�+�U2D���N���ʚ����_p��1S�"���?@{XJ��ABs�+�ݮ�����9d-�J��4����E��U��WI���2���N�]ET1�� 1H��rM�y�͂`�w��Oȓ�g�����͒�wT_���ȓF�.[9���l6�Vdus(�r��٧m~*ț�n��B�}pǎ�D{'TV�`��9�i��iK�v=�G�I��E,za_3�Օ�!�/LE�@�S�ܪS��J�z~��d:�,��������ԣ
}��qe��ţ�B
�*���3=�{�>)�$�if� �}��*K�(�H7rŤ�Nf��jg��KFE���Ht��~h<A���Sg�W�'�W��yLy
RUVH�W��Id�`��.rϥ�T��nֈ�2E�8������@��hѮ%M-3�lf��	&z�g&0�t��X�\ȩ\�.�q�d{l��GjxC���u���+�����rU�A��8`����~��;���"������������������;�%=q�)�ڐ^9�܌ʤ��~O�!������Nei]��y��딯o�S�?�k��3�do�åbO���Ӟ�$�`���ݗ��Xt�>�	Ȅڕ���'��+A`�EV�����z{��Lu�Χڌy���x��0o������d��?,�˜ ?D
��z��5�~R���������2¯*�����x-�K0�T�w�Ĝ�)1~�{;��\OEN����o�b�>��c-�� ��05��J��ZN��B����d=� `oT3͞9l��(�����`�uL<��+�E��S��n()]����՟�/���s�4�v���c��"|�cj?q�Ȟ���y�(�F�ǵR��_59�,�ѓY�F�#s޼�c���Jx���[A:tSC���,r�1�:r����*���4�~j���x��Q���jg�����(�B!I%t9,N�$޸0p~hye�p#�����T/�ܹ�lA�f�g�CM����{�6�*&kt�9MM 4��F�i������-1�NR,�3�9�sFȱ/���(7�Rk�)c��-�;��P3�g�	�aD�7a��g���K�y{��M�T��C(m�ߞ[�]����=���J�E�?���j ��?��(j�G,|Ehk�C�~��UGwJ���J@/�Ĵ��"�.�d�K�	�i��Z��xќh�Z�`m[؝��{��S�Έ6��\͔۾���6^z����~ML��]�3B�w-��P���*��7`��IQ&,���dXB�hm�թ���^M�&���p��V�)���.�[�)���q��?nT�Q}3@|)���9>6V���	�k_y˥	���H;�0�m����&v�j:5 �p���OV&p�lT�wG?M�g�B�j/gg5���}�ڏ�3��ɫ�L/�e�X2D�������xj ��@���������$i�r�2������gl���7r��2HK��GA[N ��9s[�Q[꾮r��
��O�����UGΒ7��J!��IH��<���Ig� e2}���PF��[����>�Xi4CA.;I$��)3H��sT����8� ���3C�@%s�g�}�g�"^`��w|��!�f�8��
�pE�^����-���F��eY���]������"����_5;�dS���,� �F`�#q���Ǝr�_��j��c���������N�o��7U�ˁ����]�?0qE�d4�v�qTA��#x}jr'��pӹA�H�}�X@�]R�?��'5y!@��[���A�JVf4%��`L��D�{U�ł�?�� +��-Fq���q�\9�=�`B�'�i�,Z]��=�p�Ѵ��e���fC�B�š�InNj�-i�E�Ur#n������1X�+�5`����� ��vʂst��z6��)�w�g�e73K���M��י��>����"������]��5�;��O&���b���
���Lު����qC9(�U7�aU�����<��&ۿ6@���TˤvvA��?o���96aZC&D�)G���^�!��v=џc�����;BMa,��/�=xy��f�A���'�6Z�%-�"����a�ѡQ!iҙ�fS���H~�l���B:s4i����V�T��C��8��@�����2�����q��e%"o�'��:�%��}��QqyJ�Q�v��LwԺ�F�H��V���ݍ�J�s��&��E>��t�I�J�4y��=w�����S�*o��P��;�\��EQ\@wڋcD3��{T��դc�B�V�d���ߝ�Ȣ� �\��-����s�d��Eq%7U
��%d����z�W_w��� �2�$�D�J\=(� )����1/rl}m��ds���8�,�D8�^���A�2?�;�*�\�`�$Ο�_�L�c%4`�9*Tw'�˦��]�<)��V��x��4�_��J�q$ΐE͉�x�J�R�����QԬ-]+;K4e{�O3�w%��������x[��i����&���/N'P<[J�`0��z��8�����UY���Sz�:p�����ؽP3�_�5�@�� j+���~����. �!nע�h�̢8:ޚ�6v���Z/(�#vf���%�9��8X�8ܣT��Q�^g@�H�����%�{Aվ�|s0��V/ke�6[�����5UP�xM e�{�xf���y8貯�.H�rڕ�}���T�
����)�?]6�I��,�]#V�,Y�#����b~6������ބH#WJ�LT�^�qY�g��(a�Q��9�y�H����}�����H�Sv��c��LxzB��|���LtK�b�1^ Q�´��K=Z�����2�ɖ���1�"����~�+��v3��=:T��i���
?�4��1����N�S+��BU�?(/F�c��l�
|�D�3���X�}}���-vz�����-27�m�$[��!��,���JL�ܲWk��.�� ��r���M.*B�O8���x��e#nT���;���gi�|�o�9�̭'�yM������1GZIAG*,X����Z��FN����&�n�oT�t7�s���A�����W��ʽ M{�Uƾ�.�u�@��l�M�r���&8�ʎ�i���?'G>n�B(��Ju΄�aj��1U�� �%�YY�7�$����$�ɇ�[b�rG:�����
E<�Zx��ٿv�j�]G�y�KE�մm/��š7�;Q���3O�ͷ�e�Ֆ�����(lF�?�,f�
gz7{x�B3ݕY?�N����h��B�ŤȘ>Em�.�\D:�~��@�h���nh˪�E�L��&5퀴���\0��c�(�� �qfA*Ƹ)�Mp��$B�޶?��<]��0�`�+�*mL�X�}2�kXHf
�2�~T�Y�\�aW��O/�ϱ-����&�����
�N�4ǖ?�v8z�Iy�0��9&�y�<�@	?mgS�f���P}t�>A�
�Sn�`q�=֐�ַ^6��d��O�qه��!�m(~��*��D�3��k�S�
:�Pv/���x��k�C��[���t_�4��4��ifó�'�Er�8X1�ظ�u0-����=�ǟ����oS#�@t0�^~
�y�bw���pYa��v�b��yO��T��M��eټ�ȝB�_��
��Ht�e��8��jp_���4���u"���y�H�M����M��pĕHdGQ��\�=릀���c:p1�̺�~�F[4�޿�=��K��J��o��?D�]�o7C�)��e���(*��˓O԰K&�|lA��k0�V-w��]�~\՜�A��>;2�˨������)�?���/^:�:�-�L��:#B�������Z���c�`�=�u
sW�4���-z��X<�=��F��������=eJ����E��e6�^�J�[�\,Љ��g�f7ȵ�-R�u�#�R@���}�����U�?���Ɯ��^+��@��`~�St ��� �%v�JR,�@��yd�������&�\��D
�rt�R(O�V�-��+���\2`�����%�ɘ�i�w@rQ\?�J�������b��z�������)Z1^X��p�6i���d���l�f]`=J���� ���5P�O�.c/���!v"���L7���z;����h+@������/m���#m�LW}ɓ?O�4�e��)�W~�f���	��J�6#���m��͸��H�<�cg/�G�`���6ӹ$�ʡ�ӘKx߲�V�3�#�j�~�h�wŋ\W�����	�$g�J�xx�MX�4w��_�fG�4�iP:3�/���+9${"~�dP��?����$1�ژ�|-d�5"���|tF�sc�C�9��i���o��7Q6O�����˼��T�y�1E��AAqNf���s�-���b�d|n���p��A��5��ن`����|7�=4�Iyc;ӿϙ��Kh0��-�w�#F,�DFb]��.^�"��A|C�n��+���<~%[e\J�l��T�,7k5��� Sk�՗b�$'���jFK�!V3�ч@ɍQa&#���h���_�I��O�
�1�7'_"�6(�Mq�����2S3�D	]��0O�Io4`���~;�Y�Ȇ��Y)0���{�lB�h���e����ḾN�3.I��0�V=��.Xd~۾ۨ�&� �B"!k4�}Ъ{e4�M>�2�du�vvR�����=��'�،'_��Ő����"��`�Z|��l��������@?d������Z����������j���T��,�������]��+5�
-�FO��5�t�azx�wT�����X	#��=����-h�F¾�`�]�*��D#�'����	�95$T6*n�9AJ:�Y��I �>���x�KW�7�8� �xU��"�v�����4���4)�{���[~c�Q}wD骊��h�B�A*�������ؓ��\���a�#2�4Vud� >����i�5P�\s��ypQZ�6��.��	Kd)vI�7���cx�� `�pKZ�c�wR�߾��/�Y��JRX���([�"M�e-��x\(6���\�>�uH�i�D6�e�ތ�i���i@>��UL�?�IQG������G�
���(�NF� %��7�#uJ,�L�6�J^�؈�:ٷ}P��/P���xE.�n����~Gc��앝�x�����y��)v2%���9�t�`�8�$�ba9}��h��e�88����� B�����dd���LpW����k��SuPQ��ı \�i�'>̘t��)3�ۅ�cp���G$�lpY���|�1���;%tВ�P|���|�Tb)���{qW� �s�9F%��}�`��S�=�hmmf.,s>�ͱ�ӭ@����?[�թH=[a=�([���ަ��֐���cIp� ��E
�-_s��BS�א���;j?��Z�k�N`w{Q��|b�ʌ��RH4mmD-�+�h�1f�?B�a�pH����k��ى�E>�V U��9�UQPn�0�"9.��r	[M|��
�r!i%5e^���`��a]E�>���aՑ4�5`("e���c�� j|EY�lј�Ūf���Y��.����(�����z&�G�_�ۭZzD��3�b������`�;6��OT�2L��i/k�����5G���-�US L�Dr��o��LCUR%��X9S�:w����t�-��#��Y?0g�K��+.hx�>�~%ޞH�~��a��fl���a:�����i�"G�����vGxB;�L�zV�h�w��:��an����4}��h,��+�#dX�с���'l���$g�qd�M�D=�(�t����)�* }7�\��O�-�N���E|�i{�֒}�d�Y>m���uD�Y����vH�>���ѱe%��ԁ8����8 ���A1\��w����-�}u${4�o�" �Ѫ5-��Gϯ[nbQH�u�a+��HYm%���?|����*g�R}������K6>�!ڃ��M����~�f��6��S%���IԷ���)-�T�+�dv:{$cT�a��b�0*���)@�O���zJ���i&{�0&�ω���YC)ˣb7r&�f�'������LTr��搴%S�5,�UpXLxl�*��YM���f�p�p�S�y%��+B̂k6aHw��A��Ŋnu��>pR�ug>�	Ft����f���Ԇ ��?��?%�.��.��B*ذ]H���-�q��m�bz]o�5�����Q��fC9$m������bJ=U��"��BѮ�h�`�LM2t��$v�����ctň�B���Z�P�GG8'ٶ�<�����3J���MT�)�7�ڽp�=G_�ݠ&mH�V���	��`�hJ�c�ob�#��}M3�W�D��$M����g%�㰲`�t n����3+���(�ʕ3�0u�/~�$" �A��d�C�YQ{�٩V�hFv>w(���W�J���G�v��r�C��hEhPI`%�R<� 6���ѻ.P��I�5�V�-�An1£ez��7��|�Q[��F���+��ٞ�JS�,��*�n0x�㬷�vt�,5ͬ{�^��U��ä���Y�uw��,;J~U\�7��
����k�5Ϛ؆[
pyrR:����>��W`oB9�*+7{�h�W6��������P�vr�I��>ge�ċ�a�@@��E(1���6���;w$l��&׬�7
h�T?)��v�\��i����zZV�tUg# ���P��{�3*�r2��A�(��l��E9�ec۱��}�Ey$��N�!?#�Τ��8�w�=�dvI��-�5�i�	k$�r�%�T����<8�5�$�����3�F�_�*Ez5Pσ.��~*"jNjW�Rt
�Bj�2$K���W�[��O�烡�k3���$�n4�L֜+��_@ ��$��'�@�mvۥq5�Sl��V�y7��˾X��F�����n]z�p6��d|�b@o��Ը������?�a�٘DF�3'��{�|B�93�t��E��u^��xg�[�"��'�~�w3��BSHL�W�'�f�����5��}�u�Ή��O�t3��D��BPper�q/K�8܇̣ գ/�\,*�]@b���t$��}M�"�`�#oҍ����zѳ0E�F����RbQ¤��(p.�/?Y�YC�[�S�O����^� k1��9��ρ��9��c N�{��R{̔����e�����WGp��v�}�Myg�)�U9~�O4 ;��q��%v�e��f/�����N��	u͍�� ������Geb=a]���H�!A�O���ܙ?-(4�)�A"â�l��B=sb G�6<b\��Ӎ}4��:�vV��}"���fM
���P.Y�t:T!����}���˝�0� ��5�ߦa-�K�$�n5+� �z�����?n�*�ӽJRV��@�Nh�2%���3�L`(�P�n�$1�9h��Y$/�W����gxG>MҜ&{�m ���u�F��~��;�0>��+��	���/�Ǒ�ר<M'8k)����|�m��d;B���f0�ıSN�#���{A5'���S�r��Ė���p�B��mR�=�:Υ���~!`Z���������5�%�n�]�~�Gb�G�����I�Aƅk�]<$8�7u������n)X@���8$���ij�L�/�hcJ
�(&=�0*'���L�-�)�d�������?��5�t�?����P� Θ �xߪ��������p���vv��j1]Ar������0��ۧ�Q�Ǩ8<S-4�7�M�|Ƒ�ہ�)�M>�A�Y��핓#�2�<$��w��|�JbPa�	���ū`����Y.��w����[)�Fo�Dɋ����
�L�(�l1����Y�B:���Z�sE0h��<ד"�V	..��NO��H�^�Vş�c�������t6³RzkJ���1�Ϧ'�.���{D�O��d�J�a�P��jK�}k�ix|d��$����9YK��Z�~�&���4-q���:�>?��ש�-
�!	`�ւpR4����.��І���!�
�:ȓ����$��X�FT/���&	�<��Ly���8�\�����j�b����!� �$��.�t>������ ��8{ݽs��A�ͬ�j�ȴw����·�ю˩�QV-�:��8T7�^a� &�M���sCw|m4�.�?'դ"Wk#�ݦޟM`a��Q�E�lh�1��N<��)�K_��=b~��>��l;�J�#���&���#Q	Y�B$���(v��6u�B�7�	��s�Ӳ��� �&ZQ�_Ut�'�\Q'ƏZ��8�t�(�FW�AI�I��%e&��ӬuB Z��
��]�>pZ���H3[�&J5YA�o��i�4\k	�[y5�.ƺΓ6ګh��!o~��n�r�>�:�A��pB{��i,���@C-��c�sf��QheI�J8��1K�����~Mb�/}�����_�ο�OkkDi	��mXn���YМ��?�>������Z��=�0�2���r*�'MF�O:��B���_���湩B�|���t���-��}Β���D����I��Y����(����e�5���#����E�8'�?0wB���b�6���x0����5��
�T���grA��%x5"x�d�{0Tަ����V�$�8���u�e�h�� 1�
mZ��(OW�u���5����Å	��:h�@�m�ĝ���rQH��%#:�b!�^=Yq�7[��"Z��0G�c@g0�a��v�d�w��Ϊ�:؞7�3��Pz��u��L���~�� \v8�Ƭ�wR�>͊F��qHq_"Z�q��<�<��A�	��j!��^�����m���h&�|q��W���c|��K�$x��4�k�������J�!p뭲?�(�ǅ�%!�rV�B��`5zR+��1w|W�tD�K��n��%�;�� �HP�<Np�ME�#=��U�&B����i-��Ǫ��t�>e	���;�uT��Էc�;}.����e���}c������0`�[bl��� 1�k ��	}Aӟ�d��S�9����+�ڝ�M+�>�e[�����l�IO�F�jД|�}$�ݲ�Q�C*ǽdy�v�|56����#z)�V�X4q<��ޗRڳ���H��~�N��_��9�#�{�j�N4iR���������N�Ԅ��'�;|���| wF����?cϥH¢�2(���$�/X�J��r��K��vm^n�ܪ
���"�û#5Ǟ�V)��g��!��~W�F��W	���kw=��fe� �_Y|cvV�7��Z�z�!F��Mۋ�ҽj��Kb�g2|}\b��Jk��vR��L�1�*R�g�,���:�<#H���p��;�x�F��B��u%�%濲eI<�j}[���+��.1��$G7#�ئ%��l���:Q.5�j��S��u�Ek^g��m��(r�"W��hg��������!����H����gl�)T����2q��Ȉ#0�9�T4N!� �d?~�s�"���(n�9"8u=�u�PîIaO
�7�G
{�)�����F:>��[���H�%w�`! K<��'�2�p-	��l��$y��gG�Tg=t[�靤I�
�L�\�!��2��uwt�m+]U�K����bO��F?��^?y �R�����S�i���C`da{�����{��0\>��1۽$��[��&��Ƙ�A>�i�W��f�c�F�uTX^O� g�@�ydڭcX�LzI�=@�5R�j�7�QK� h3�Ҁ8���K�^��$P�np$j�+�m�?�y�P=ki���:�T�F������,%�G���a�I2{�l`�t�=JՉ�а��6{"�Μ,&%��N�=/]�^���7��ω��j���&�'f���	u���Z/��ٷ�8��H굅�f0�0��&��u�ﾡ�5}0'��S{�$'����[�ʑ�h��M�@3gz�N����0���sA��:���	VS�n��|?���	z��C��Hr[�wY4o�G�y�~�9w8C���r#�=j����T4~XV�������
��JT��C6�{ǐEM8�
L�V%]��WV�����ԙPF�:;����0�V�����5�0,��<Q./�x=������n V����;frV="O��1�9:���#!���"C����QN!q�pg�π�a��xH��{�Uԟ)�.�>��p�|�Am�"��e��Ll���^�D�mD5������O��D�X����(%��p���ｺ	>�d��"�m�\`��?Z��8�ƶ#Y�#a���͉��B�H�.U��m�E�"��
�KC.t����+���.I54:�	m䳙l�7�d-���4�Ɵ�Ib7HQ��G�܃g�z�)�~-O(�h�$I������ıj�z�7��!��E��lpX�ȑԙt�uN��b!�=�i"�&,�!����6#�\�",�B��Ck!�N-�a>q�n��D�x�C�*>*B��X���;"�ڿ�#Vٓ6'���^ek���=�n��k��C�J������v��N�cwҍ�J��w�\J���w5S7��z�ʿI@�N4,X��d�+��ovS�=��F�E���j*�s�*���ra��f$�������Q?J����"�Y�Ԇ"o�Z}�M4����(�:�a\��bt�G�UenCk�K�a�#��D&�^ݠ��U��ɡ�V'�x��2����5���]��)�Q*B��#N�a0�#��	�HJJ����E��'�����=�ю%f�w���;�T����OA�Z�qo�
�,s�O��M!Mv�\Ξ�t���� k<�&�p��_�_q��m��C�������һOA&'iw����?��i��FB��͹��AK�&���[���I��'�h�5�	�� 7pN!�,Sc�D��#ӿڊ�����}N�A ����������4ÎSB6�5��q��x�!���Y)�1e� fs&��B*=^g�&�+�QN'��gT��)�5S)FX�O-u�u���44���״�(�7v���un�v��*2���M��bTLes�m ?�>r���v	4�&�@��Y �f�{���6x~B���[��>����v]��Y�vN=�M)���$�������{H�u��ܵC�|OQSҏ�ٺ����S��}��옊FO:���;a��@�n8����F�j�X��iݢh�2�i����޶�����r!ԛ��RWf&%���NT�������XQX�����'�'F-�mV�r����o�z:��T��V��"���(0{��]h��~�#���`���m�`
6�@�|}�-��g��@�!bP��� �cf.����(�x\\�[���U+,��B߶QZ�͗��[�����W��b�.� ��x�߇U#QLe�C�S�Z�n�T&��J�@~�Y�����9o�(R琅�'��6[k�B�/R����a�c�+�@@���'����+"L�n!�bn�AϭK/gʗ'��T����_���U��yj�D�T�9����fB#%n�Q��jk��`�����!Df�c�;3�u�J��#xW����&l�G��iz�3�y�F΄�xu��$�tt]@%P�XN��e	�h� 3�֑8�js)��п�� z��w�W�/iܣvܒ�Z@�4H��v1�A��`op�-�3�JHlX(r��Lb ��̦�1Gg����]��b�H����힣����m'$��T,��lg�|�j�O�*�3��0	3��%��v`)�Wi�����浉�!�HGR�Ms�%�ޢN8X';Ƴ Ր��*ͱ�Nc�VH���|��Nn"G��=���;���!y��!.�8�v|ք!K�Y@��:�c��Pɟ��*���U� g� �Й��Q&x'R���-C��vr=X�|;>ڼ��	=��	��=�Q[U���f����c$<g2k$J�5����/�(�\R͓"�shה4���CD� �����=~���c9���vM�P5Q�g�5K�J�����C������!(���}� Y�H"�>�iWP�%���Fb�re~��