��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&��n?��1ů��> K�-� �&�T�Ek/ֆ�\�놭5�DꢘP���+L+X�4��J��#�0�8���������l��jT��+�(���������6�MC!D�;�m�퓊D@v_p��䙋ⲝ��C_�6�Ռ��#�� ���	RD�4D��畓7���vn�H���0���fX����4 �CS�C`{��;�L����li��� y+����FD�p"��]���y��R��K�({� .؜M�������	^5���ɋ��&���&�@*���
e�� �t+���
_6��O<��7f�M��u���m(MrN����z�jL���@T`��M3��c�uQ�Y���%�dD���,�~^���y@Ga��(����C����	��G�86�S$��ɳT�ز8���:r��/y�[ݦڍ#A�����i�&<nU��<[5)�Z�-Ĭv���0t���d���"_���:�'-��d��*��q����_d�y�N-��~";#��������Y��؆���	6ZJnԷW��έ$Y�K�?�4���L�w�Wmiɶ��Y�?jx#*�i���F�m�E����O6T>]i�_�9;�!(��kH7�OS��_��[-M�((��lO�s�$�g�x7`��ZV�E���F��,9�j	@���]}<�ahb5~ãdl&I^�	v����-�@�@���	��!��d��`j[Q��� r��;f�i�.�m+UH7��/OV��c��������l��i��M��*'��?���G� SK�M��H?�ç��q;��)��Rȩ�"@���r��Ml>8!�S��L��EgeH]�8��>]GR=&���C��i�Za�z�,�F��h�q��^���wT�a���%�9�n��?~SИſ~�mu�OlIv�4'sT���/a��^��9��*��G�Fh�DM�_��CN�<�_Pg��O5��}s�%��m�o߫R���X�Q?��dK�Z|:�=��y����&���O�T��<A��C�1����!"�N��4~���r�5�.��������R[�9;��u�<� 2�X��%R�� �|�ս�}:���Ey�xlִ5
���}����ln�ԟ���ƍc���3l�k�O�`��fX������n2*H�5AZA�?_.d.�8��1_O�&�gy������J#
��A�W\��H/4�d��Q2�)��!~O˛7���<Lug�����l.�UM�_��6���E)�a��!�B,�4ƛ?
ϯ�$���J�`f���]����^0�R��e�Ϊ���U٫9�~��i�%ӏ���A��U�`K�l���A�:���:�����7�CR���D2PK�B#�hx�@>>_:�����
I���B����Y#�G�:㦸�����]Pdv����؏0uJ���}v�g��������夫3!����Qc}b�ݍQ�p�^'��p�5�!��$ ��,�A6���r�r�>�e������?_i���Ȃ =e^��(�"�+�]kZ�%(�*:�$b�oMch�}'_�����O�<��@�&	w"��b�~Jk�R��ό4Kq�H2w�fhob+�+k�C�z�eR~�N���ˉ 
�2�m�ޜ�J��.G�|f�T�9��w�)�ß^��e+�kL������q�/'|�W��U�)�ľo��M���M�`�!�O��Q,BꪍS�d���(zK/��7�׊,���������T ��{4"�h=���ֈ)(�u�ݬ��؝uc�r^�g�?������J7�1��6aî��3(�{ �[y/���A'��ȸ�.Θ�!t�h���!S̡>��~{U�B�9��'z��D���"4iK ���MQVݕ����|>�������L7nt��w�p�����pE��t�zy���HY���Ppn;��4C��b]B��n����ݍt�������
��p�g��5�����W�`Uy+�_)Q��J���2\^�[�멢�f�ɨB�D�(��zB����wYgX^��V"мTM_��S���;�/�b�
3�[�4$��@Eo#/�ߓ�pS��U>TU�F�_μ��G���d����l�M՝�:]�/F�ݍ�;@��QӢ Ca�����*�o�~��CdC��ɐ��1�wt�t���5C��W����p��x�s|�,�h�E�js��)�8���@���g�,1]N�?�n�����7��m��%b�?��ڃ�7��軦�P���T!�:^�u��l�g�^�4���ge&i1� 	�.ht�9�@����+t���T#�_�լ��@���@+��ݱ�hc滦p��M�Q8|mk��y�7H�t*O��Ӯ-�͹��Эŝ�$����Q���6q��lgH�9q2�jc��[���`���hC��G���)/��饦+@q��Fv�`^$X���i�ʯ�o�۶v1���h4
����^��^O���B�aTC
�Q��VS7��Z���y쩊���X҈�Q�<!CQ�F��h�/�,��f��qvleO9�+��J�g#�^T���$�/5Ȝ^0�L���H���u[P\��޼R;���4`�׋�s���)�81�qF��ui��"���m_�_�-?�V����~-V䑃�)S�%�"�4KNr֣��$t%���ps�ul�� �X�r�ĥ,�����-��Z�"2w����!PG��WW#BY$��?;����j�:|g.,Ɠ�A�p��w ��MM8�(u*�m�88 FͶ~[�}��wR=a-�̺[g��Pn��|n���Mݧ��P��r�{5�\o��J�����뭆����UQ�T��BW���A��#7�զ����:.�k$V#)o�"*��������GN�d�tU������<E_�{��6�ľ�@G�2q�����f�F��gbpLO�k)��2��M@^�]fO���@Hn���䷢�k�	�Y3��AR�ud���G��G��S�o~�	���v�?\��7j����������wG����x��� �3����-?���h�tf?f������ ֚����|A�I˫������]�:��|[��Y�2��q^���W<<0��yz;L����������K�ޒe	�O���Ķ���N��:��q9�=t�]!��W�\[$ �ǟ�x&O���ޭ���mh�⭛١��хkx] dly���x�ǉ͆�a��3Գ`K�x�m�S4]�9�MBS�Y��trk{ew
'dA��]`����3t�Is�/u��ݳ�^a{�I6v�dM�/KN؛�ڏ!nI>�,DO�g^�Q̘_�:�X��䴧1�ךs=Ղd���-^�8���l�r�9��%�1�JZ&'Ӭ���U�N�u�}���w�ʫW5�V�O1�L��f���x�������F|���Ȇ�Z�������c�&�T'�YXz��B[MMC����ב���z������������ѷЋdb�L�HH��&��[�zk���@i���Ԅ��d5-/}����D;*�w,\$�bA�x]��fÑP�x�,؂ڭ.*���I��}�Q�V���]�n��A���G-� <%V!��f��5���.=��H%���5�j�w����Qo7ѣ�e� )���	�̳=��Kê�L�Tm�O�'eA~N$ϫ�V��1r'�mZ��0�NJ��1T �A)��b��o�M��=�Hp(s\L=�*U��)���C�?$�i�v�Q	;��$X�M/L�Ò�����:8uˠPϭ���!=��<v�6������Ru���=��@�2���߿�kOZ��9�V�/�u�Qd�
�?r\tn�%�3h����˓�%�~��0�RԾz����lc�  ��>�s���'k\Y�\�M�͋�\�L6n�CAh@��K���N�mi�
���q�X?V���ی^%#�p���O	_�_�?�q�i������{~j�󫕀�V�v�c<@�G66��;��P~t�
��|^n�SB.�o�W�]�Qqo�8^@
j�3Q]�>=��A���E�R�n�A�?��s�0F{w��܆ $�D���W%z���R �f������Nl�	y[��V!�^ا�	�I���̹d��L{���� �6$ʕDL��I�+�⑊�r�iJ۽�=62s=�c���Evv���,���#�v��1�G�����W��/�ې���i�������/%���LW?/�.�?%��:�8�#w�T5�+�[��6y����@ ��:�"�Z7C4���GH$�e��u!�lc�gEԂar�~��2��54:�0WȁN�U��.��#�C"��Ӹ/h֑�4x+���W�\���hU)����#����R�pK}ֵ=�ͫ��Q�k#�$�M��#+�Lq��-X�C����7y��ӫ����� ��`5+�R[㫧�=$�:����>�(���u�=L�uD�6��=�#��/̨�t��jq�2D.�P�&H���-�u���f���n8sd�뭓�W�_�k�l�Fq91\�v[��\��gğc�L4�N9�7���^�)��f+���IN�/Ž5֠�|'���E��̷WE-B�{]:k�OB��Oh���_�_Q��-d���X�B8��	{N���������	����g�v?��Ⱥ�{&6���P��@nI�`�������t/�N��9������#�{WK��+���I�I�X�.,�sW&�Ir�����9�,��u��Xho�ל���4 ���7:$�9�K��|�ҮN�6���6'��㿮4Ҧ�Ef>����b�	��uj��k�?7MG���ްP6�Fr��o
�~��M���^L�1"	-�ARފ���=�2�ÒbVX�;s�ԝ�9h�q���}���5ߏ��׫�&�u	l~Ց1�{�6����/��S��ʦ~q���le 0 ϱ���� E�nM/���B����q�E�M�:�oi1cy�j-��(�Z���)G UM	�`ٓ*��E���Zo${�G$N��vPU���vd��(L��~�Z�^�6_�kY\�E�~���)�E���"X9o= 0���q�\��N�*ߪsc`�F=��'���҅�������;�t1d��&::�`�c\^�N�;��ޜ�o�2](s!�h�|�0�\���)�?�u'�R�0�y��s��Ģ���e+�
c(�������e�����C&;]�����)"�ͭv�W��H7�6�\�>�(rǊiDR�M����x�<Ɯ���醮���($sc"�̓�Œ��PTb��l)A0$�
CS(�\�P#=�7���m���G�扑Jnʬ� ��؁�2�ؑ�*�t0�x�ǽ�`��߉D�U׌�;T��o��$~���ʧ5�{D�1z���Ro�+2���S. ʁ3-�*���*Jp��tb�}d.j�[Z���`��� �]Q�ؖ��irK�	�W�C#
T8�7��x�C0�܏���8�O�N�&%?#�m��kW}w���(��
��t�]�=Q�(�8[4�
<S��Z��+m�8�N0�d��$�V.�j�"���?�L|y!�$|�J�C��/�����;3�+���ڿ��*�*���$P{+!A�di�?�Wcݶ�����}�����t�'7����ws�5Qc��]7(q���1�f�U�~����$�^����p��i��B�
��n�������jXâ>?�G�m�4w��Eػ�A�֙v��( ��<Qm1LL �g<�cZ�lF��9֋�t�ٖi%������8�D�p2֚�*msב�������l�E���y���lh��ZR��]���J��a!R�)0h�����	��������7�}��^BW���̼�
n��v�{�u���V�I����Τlʦ�-m%���?4�΁��r)��/-Q��%��B���9ׯ������ڏ��6����	�E��%Uc�9I>���ky�w����)[��u��y���� �&�!�'�R�Z����ؙ����r�!g�#�������K���eXi�]��M�zU����Tl�#6Ⱦ�@��yp�$��\#xѶ� -��.�J�!���ҡ�y$2B)�> ��lLz�q�$B!�%I&f�K���~Pm���6�����J�	"d��"�R����9����(����-o��3پ��!�{&̋���e��mW��S+(��#��g3�=�(�2и[�[f#�ox�� ����3c���V���I ��v&���#@�;%kF�m-Z~G#.��:��d�#�T*��y�F�+��Z�k�Tzq��x*T�l����5 :�y���F0�Ў�i����-�졦���GRR>,�	�6C�2]�`!e+Y\��C�9�"5�݂���<�׋����Sө�/�"��O��Y��X*{���n��X���Xn딙|up��B��0�Z�ad����g����~.9����&pC��zf����F� ��M�����@J�Ӆ&}�t�!�7{Ik�I�q�o�~J�<�+F�S]�|�MF�A�{v�H�5"��n�+}嬏G:�n�J���e ៪E#r��� Z��L�6O����E ʸ��9�s$/�������y���w0��4���ϥڨ��F�պj�h��G�o�e��D�H�?�{�� ��:!s�.߰����a����˹nJ!�)��%ot���?%6h���q���xtTN����WBx�˯o�g���U\�Uձ�v�c��ۥ�R�Á~�j���c��wZ�a]���)G����b���O���j�([ kI�R9,�I���Ado#�Ӊ���a�rf�x?H�Dg���M!0���h�=��y/;l���-�њ\ߠ��2�E.ng\�8�Q��O�H]nQ��
4uBI��G8oh�7�J��cƢ��:\�c�����"�n0�a7������I�}xH��� ��%��H(JBԒ`�
�m��c�K���oަo����d����(��qaw�a%F�:ʉHA�se�yy`W�b�ˇ���~Q_qN�a�-u�A�ߔ�8��:���u-�J��_�%��e�~�_++
X&���m"�g�˒�����1���'�"?�ip�N�S��Ko�vi��)���,�P�#�B���"}H�A �l��G��P���U%�sں2���/��?t�/�d��5��ǅ�f?s0���A[a���B�Bdl��\��d�%��E��~�c�rA�Y����)�zoB�!�Z��X����Υ�'o1Q��QH��Q�NT�Tc�U�p[����L�$"�����k:�.(�Out|��~��L�pk�I�]`h��"&�u{{*�7�o��XX���"�>����z:~���w'����yg�p���ܱ�����W}N�t'�� W�yI���B{+����C��/e��޵P��� �gW�4�;ǳD^��1k�y�6�)ռ�m1 �u�6Nx�R�x}i�Ai��l�d܋�!��&�
>:�!��}��?;�WU�؃�i��!���17�h�"T����R�`����Owz��p�n����Oe�!5{[R5�c�����l�x�@:�a&��ϖp�]C�?���[�OY�i5����b߾��,�̥�'uIrDZܡLE��o6Rwc)] ��;o�
m��O٣�-c;4aʄ��#j���.۽��;����1��@-�_�i%3�G(�_G��; �z��X�ל�D��,VG	C�)���@tfv��<*��UB*w(��[�Ք�_SX{EÆ=��O�$�]g�Ρ��B�����5�H^=�i���^(s�lu�F�(:�9�*3

4�����W3�������g��?_(F3�f�����$V�;Rg�
���&#����p�;߈��p��](��$�����
fK�βaK[���~+J^�M�U���`E<�L��zs���7���E�Tj��C(v�~�c��{"�����!�m�͸ת�(��Wه�	d���x�Х�п�:����94ϭ�u�v����Ȫ���h*G3	�T ����B���;}�O�89{�i ���u���D%g�gx� �;\ݸ��_,
�V(�-���9�j���:�c�(����^����]��df��{��{�'`����vB>^$BeW0v�".��y��Tn�L�Ɵ�	�[���!RXo���@�I���F�Kk����~b����$�iI��[~�f|��IP�Ǭ�L$���41+k5���<e�#�/�k`X2F-��5)�}_z9�qu��}+�y5!�'�X?)�+��T�����ØB����9���0�n��x���(GB�Y�����jZ�	FF,s=s �|	CƄ���I9�q͋>��V��A����W�7a�����u�[�AO=1�/���>��ۃ�r��ą���@���;�|�G��U�uCV�:���i��ۖ��7�K�8�>���}�;��/��l6�D�Ȁ��:p�SǮ����GN%��n=E���C�����R>9�L|3��n��V�E���y��&`�vY��#����&�<�Μ�e�L�b"�Ru��DƖW�ͫ�ox�_{�s�w�P�#��������C�Q�)�c-;n��6�7�3�?�\���M���چj;��]Z��:�C�5jrvhy`�p���	h��װ�J�s��Q}aM+Uv6-=Iڶ��}�4�P�諆F�pt�(πk�������	��|���&4�xsu�c����.>���E{�?�x�,����F7bj�<Q��h.]��̪��ס,�%>�}~$R4'�(�{��'��
������A~�8�M�����P�-Y!��kp��d�aC��B�s�"���4_^9�#t����^c�//��3����iBB�Ī���`��[t�G�F'n����)���y���@��r �{�r�YnR�Uv�l�IQT�@#��/&���]Ċv����ĕ�:;�=�&�Y?Qe}��56�6�[���<�YVn=!1��F2`�.������E�iT��b�q<����gC%��/Yɥ��@*����u�y'��L���y��c������"��o�` �i�a��0v�GQ�dM4��Q�/�D�#��RV�>�s�΃ۘ�����ؑ�͛�Q%7�K�kӠ����P����H��4���� <@��>�f-��'��kXY{�an�� �YY����3����W�sE�A�e�GW�!J���1� �Ҹ��+�����:
��[����mn�рX����4�DjK��o�I�B��^l�yiCC�C�����ԗ�}c�V���������Ci3Bo̩"���ɪ��w9HF~�}�p��
���{���+��ѻ��q�Y\��M� Q����E���a
ډ��
�I�ˑ�b~�Ϲ1QQYz�^�2��W��Δ&n`�?\�+�EO�n[��oE�F!G�JQ�����
9|���16����^As�݉�j�d�;t��ˤ�r}��P!ZY� ��@�u�5V�PN����2[�[�q��zr�a9�_�������� P�;�kO4K���t�<�5M�D+d�p,ې�ܲ".���w ��!bo��\M+�@���]#�j89�f&I�4����u�iBjK�d�8�b��fQU �hߗz�L�!%B;/���1��q]Yc2ag��dz8��7�}y�sQ]�n�a��E��@~�b֮yꔣ��]?j�VK�^$s����oH��	��1I���d����rk���.������K��`f��.	D�/��f�u�� ���Ӆ�ɏA���J!�H>��溞�^a�>�C=+�w�*_ȏ��_�qWA�M���� �S�Md�xr�~g7�Tz&~p��:�x���:\�c�^?ny	����􅩡�P���ߩ�tu1/�r���P����g&�<�!�����4c��s��?��1)
���5	gU=3f�:5&���&{�'|�����o�'X���e���?6��Ʊ��4����|ms�������!>���ҋS8z*e)��=2A����P��Γ�����V}nAA^38����%Iج�z����n�d���i�S��Z���2c/~6ڐrN̸�D:����(Ig�Z��َ��%��=P�fPc+��|���d��WG>1�ML���T�/���<c�E�{nʟ���s�NƑ$ �.�s~¨��\��Y)gE�PE�;�}�v °�nU$��C�p�]��D�4�� J���#�>��;/j�52�.���*�=6�8k�������_S����p�`:=�߰�y��M)d:̈́;`����(ug��%��#Ї8�7���CU7�s���f+H��{�*�rq����7H��d�s1��{<B��$M�����Z���I�^�̰�es�H^("F���,����}bK�r�aE�tMɨ%Rn-�V@š���e_������ܐ$d�?2K����f3>���g�q�ڊ�w���z���/�U�T���E��"����8NBmB��^,9�~���#��<���g�7�P(�"��<�{���0
4�=��bO����	�aU�T|�ˢ����(���xG6��\�� 3y��M�Г2 �N�͜-υt�ѻ�Y)����P�'>T���n��ݹ2�-�a��p�����u0q�~�v���/=를 U��!:+�+���^��,<�q��9M���Uz���M�z�J |yoK�D���_�����c\:��u)�c�ʀ�����!Y��@�\P�����bxb�wB>e���v�#\�hn{� HJɖf��v:��=׹x��M����//�	�lM�B�:��I�'��f���fk��c�W@��a�C���!��}
bZ�q��F/�8l���h>57�H��x uF��d�j���1n����o�:���k5�"����j��|R�!��m=����ۓ�C�[v!��8�0�Lf��;\cf�g1 7}�id�7`0����߷U��o ���C�g��M�=����̘�0x~Gl 贅��P����3ʐ���2D��񙂸[�p@Tï�\�6��9��0��Rz��3�^��b����T!+X?	)VK�|�·�AX
l�u��h��}٦J+D���"�	�%���ÚڎU;����61�ƈv�l���1s�[�	~���}�F����Ǭ��Р'���N����@�A��1���I��V�h�\d3����Oh�[�6z��9�P��Y��T���z*�i�	�^�W.|�|�
������~E�w��]�Y�қ֚��\7qO�.FO��Eĉ��G	�A��
=J��3�bm:�4�}:��Nl�-5��X:�-\��>vX���ގ���L�&�1*����3&9o���Va^�XA� s���_��$r!!��
<9�cd���H���	2.���w��@bqS�(�V���dJ������t�3�|/���>�? �D����$e����g�N'�W�i��
�M�a�;y��V�%�e%�V���b�z��r��J�>$a$�r֍WoJ�0����5Vr|Cfdi���u��.nV>������9+5-�Nb�nT�DY��F.��0�N1�GHX���	����vgYAu�}2݂'��^^����O�	>t��4?�$$�߯����S��ojܛͱ�^}���д����G�
v��,�n����3�!�h��N����T���,�!q�&h�h> *���TQ������k�`8b��I[��J���V�y�e
Q�->h�o��S�-ّtj; >�5�vf�� �j2�Ig��m,N�W��P�`���.ujM����-��B�==����b�3"�ȹ���o��"�跚�����<����?��$����}�$ٚT[Ρ�¿%�%��u�!�4ڹ�C-��m�xF�d�ZA5�5�Q��H��r�b�~1�	�������G}GD��z��뭈�^y��Q�<Ppl���J�ƣ��l�-��.�_9�)1/H]�� ~���{^���h����H沝�U���P(���V�ה�EM�C͕N��u�[��q����s",(wA�k�E���ҧa[ ���e�j�����eg¨yA"~�����e�'`y7�u���< 1bo =E�,i�������+�-��L�����8|Zi�ƣ�<��^5o/���E���Lπ�:2���L��e_��ݱ�ٴ�B�n�l�j���'",�3�,�5���R�'�E~Z�
���sŶ�k�g����QWŸu/�t���7��A���̙�/A����|I6���m�\\��b�NA�-���A�zٞ�5C���`����,v�Ӡ�vu 4W$i�A.�Y��L����2�q�I�'����f����r��#��j\	pЌ�p�Q�02�f�=�n��
��	�3�\F�v�:U��a#�Ϡ��IEKF�E�������Eh��%�*�Y[P�q�&���&M��@�&��Zh����WtQ0�rД]&�H,�3�]ߨ�̜�ƠyD�*���K@����k�%̸qYv�sqa��-��]�S��H��|%@O�%0�I�2���L�T�p��9�G�
��:��+X�Vx~��wh�����;8�}��D_H�������w�P��(/�̝�)/mK']�XSk�g�J�q�֑�f��5C�ܲ?�4r>��h6�U"�`3�f�v�G�JC#uP�r9T��&��UmZ�k����+�c	(��C�]G�v��zL@vo֢A5�ܠuN�ў�����P��������_%1�U�*g�������15U�N�m�,B�ȉG�z�H��~
��o�ʛ�A��:�{��|$��]]8�B-��<��?NG��H�F8))
]�le��/~�B2"lZn���'z��r�@g��kky��h���Yj�]��U�4�!t}a�1�c�i~n$�N�7����@_��Ϡ�9DXv�RySK����x���5pƿ��f=zs��F�)'q�>���uV���������/ϩ珝3VC��P���|���׮����SG�S�=B۶�� ^�]o_�$��F�1oAە)��Hqa!�� 2ZU{����S�l���;��b�K�2z�d`ɛ�=���K�X�@ˠzWS�R�,�#��F��Pe+M�ex$F1������MD<�ua���G�҉��\�d��@�`6M��6�����X�k2�Ⓠ�}��!P̍��"������]���*��ЇWOԟ?в\��wb:[ҟ�f�z����q�k�Ӯ���#I��z�L�#n�lo?�ɐe���ZZ�k����s~���,��&r4U#��7�Sܭɞ��69o�����x�p���]��v�W�ᥘ�[N��-����Ȟ���3Y�6#Q���z��P��[Y�N�2U�(��*��L��́+{d]�'O���-�o6xlW�vs��,�K�#���rt�k�3$c�"�3�B�cf%�m{��4���|F�Yf�n�y���CLe3�c�K;�|��MU��4����K��a��{��61��6����@!|�\<Ϭ���ѓ���� �!�Y��mRh�"�m�0e�zD��N�@z��S�$8k.3��V��>�&oph��sF�ݡ��X0���$Xg ��ϐ�[2/����ߕ�;��R���PY�!��||����73!���"�QB�K��y��=7��+��7�&I�����Q���6V���t�(Q��uM�(��<�#�}��l�Ďu�����G�s;��)��ݲ��J-�"�hq��f�#�J���2�y����ГշOf�gJ�^Y�"���nN�PBʌh��7����E����d�䒘��ȭ����ݟaU����G*��4�c�6a�Z�9YSۆ�������tn�[�ߜ,?����駢?��(���΁Z-��[i�S}�'>e��g�����W�pl��2����]�e��\�V����L(RP�GB���,����d���!c��AMo"���N"	k�h���iWg�q	o�d;�K� �'�|S.�0��X���f�0ħ:G�T�PK6��'�B��g�$چxK�#�	'`>�X�58W5�.�@O{�gX�@?Ҝ��kSzt�Y�xS)ٵ]�nrauAc�2��9���ī_V&l6l�����Y��B+(e�Dy"�Q��׀Y/�0�e�H��n��Uv�&x~�Ls���{j���T5p7菰�ؗ�$��ľ��R���9Q��4I�(U{����<4�W�x�J���yy�C��6���h�_�;}�V˰7|�`rcuŔ(��>tc[��*�{d%��4FO�C��O̍Oc섷�&ڻ�$S�p ]⊤m�\H��? ��H.]Q�������W�8D�6(�߮�3/�գ�b� �W��fR���LcS+ƪ�������̃zZ�y�uď;�s|��i��7c�ī�C�$�h�z,4�U\w0��8o+k7���c)�si�Z�~�y>zy~�s�g}9�򟐜�XN��QA�~�}�u��;�E�	ӗ����ԫ�+����{��8����0�rm�pk\��z�~j���{���=RL��g(���Gl�3��H(���D��L��f�������d��ûݗ������48g��D���h�/�H㨆�9hI&]��?-Ӣ�4��^���$����yq���2�#�g|��ڐ{ѭ�]ɭs�]I{A��LV]��Z�`6�5ԍ�
��|�ӵqft���v����7R�cǗ�>}�8��������T��zEK��EW��jE4�R��?a��~��<$��cɲ��RY�yl��_���� ���/�#�'�a}i3��C ;|_�~FLx9!�4u�Vk`c� +��P�D�$�B/D��GC�� ��7_+暫��کI�QuVQ�&7���r�n�	+]W��b��%d�d�0��Հ(y�4�(7y"��w9ȫ,���y]G�������vV�����1e�no�.�{�U����� ���k�6eTSpg���*I7r^��f`�� H��{`'LI�H�u)�/L(��d��c���o
	���!@<� �fp`��]U|ԡ�t%���v����K�+!��:EK��Yb�Dэ��t
 R�E��N1��ʱq�"h�Vm��NJ.�䴀�F����|5�$5|��)!�n�uB��kQ	c�F��W�&DRbg��)��n��ߨ�A�:F�+ֵ~���8��O�qu�a�Z��8-17P����[�E��hNǨ�n�cF�R����^�<�HOCT&BE�BG���Ӆ�����պ���i�q��o��3�'x�H1�*\�� A3�e�;	aI�c<��U����B��Rܙ��#Å�@U�I86|�І����ٍ���ʙRڂ��/q�t�����2���U�p���
`+��zB����L�E�&֓�&G��"�b�@lf������[�a�)��B�T�H���'����f�����؝�IN�ě8���]q�}g�m]gv�p�PKi6N��s4�'pJsK�n���З����؟л�7�1
8�p�1����.�l淌z�B�x�O�q4�}�1u���8~�f�mB�w� ��e�LD�.}"j��b�!�3�s���y_-W�le���W��&<���)ij<]F�]�^N�Ns�K@4�<RL�S��� U���6E�����Q�f�x�#Z�O8�.SJ�Y�2��A�f\WJ�o�����0����g�D�[�.t#��vq$V �Q΍2�����1 ����/W;�D"�m[9'K�s,or~�S/A���ku� ���>~��	����Q-.+vH�6#�w�b�1'|��+��c�=�����N�]���?aA~]N
 �ΈK��/*� ����`���L��V�����Ur`V��y�jfj�v���F����⎆yK��<{L|��eU����ԓ�+U-~܃5ڙ�}�%@F�d����c�E:T�O�c,�8��AK"��B��g�ht����l���/��d�����'�,]�}*�c�Tz./���xr�D!��<HMg��^h��g���?R$��eV|I��dϑDsF�z�`��Cpbq�(�%2~b�48������S�����{�)�/%6>	B[|/^����g7�����x@�8��.~
��@���dc�n��~���k�|\��)H��I��,a�G��#����e}�R�`�����,"5�=�J}P�BF�'��}�q6��=��� &A�&%Bb�����d���/
d��M{ B������k�𦻋6I����c˯(��/!���l���i�n@�s�����,�:rCڭ�%4!Ȑ3iZ\����6Rn~ �i��ʢ����6h�u�r����ϫ	f�m1ኹ)�����|:�P�[�.Dn\�&�l�������V���!�4���B��ٸ�Yl~Nf=��X��>i���v�5EP�$m�i���h���F��k|9�M\�u����9\=�u��%�W�6Y8[e�ߢǄ�rF 닅����c��N�.2,Vҥ&�[���Y�L/Y�a�٘w�B�Gc"���B;�$�PGNrR��ȵ9 '��ǰQ���\	�ZI��_���#���n�]g:�E'�%����
g��FpP�$b�tKA�����������D��0��~�`�Mp23�.F���F���O�q�W����2��u���#F8�P$WS�(R��j��1���1��l�|�a1.���Ƨ��kV����a*_`��f���$�l�d�O��6�:TB��&������S	=��q�%�iC�|2g��_�^?���Ļ��s��&;�-�s����߻�l¸va���o�Bҵ�ԞwEky�s��1?;��a�3"f�mY�����~M%�wr�64�
_�tq8[��6��zN��n%��\�a �p�XX��ؓ����LCٯ���DB���%X��f?X�(
6Z��:������/�9 �g�?����K��m����+B���T�H�7)�O�T;��76�9[IscǕ�i�v�P�,�&��i׫����<4��w!4�-^�5Q�<���oLpT�\IT�A�7t��K�ZO؁t �}H��|�;����/`�TN�K)����)FxQ8��5
h'L\Tx��v΃�?��U��ȱ�U��:@�}�?~\ԋ�q���oH�@#�D��Vqz��)����N�D]!�x|[���*���Q_�U��ȧ�]1��,�ިd�h���;����+u�e��)Y!�%CU��$Y����~U��z�ׇ3�TG
[�s;��f�ꢻcw߆:P����T��U�+�r#/� �U�6;�Fά0n�±\�Ukt,7glj#�	q�Sae��RI{3�!���0hv�&S��Kj¯x{����.��-ۿ��:�:�%�7���G=�P~38~�_��K��<�#ijP��k�S���	��PB�����`��{�����?+�GB����#����=b�dí˲s�zS��+��AB�4���Mj�`=4YVg�+᳻F���b_�z�v��F]��˛n�#���hSJ�_�$:���uY��t�*�ܱ`��c�q�c4ݝ��oO��b���5<�ۤ�F�=��|�Z��n�����������/:��V�z�G� N�4�h4W!0��Lg���"���?4�iy���n�QT�q>���H�Ҧ�4窍�{�����ŵID֘�<�7��:����Z  ��ѦƄ�����'�� ��ش�$66��F�������%oOB��S�����6��m ��{�V�V��s7(`�K��]�[��!e���PR@_��'x�A��+�oz��u�O�o'5����Ҹ��	"�Z_9��d0�]����3}� �ԇ@^�Ǐ���sl��֟�*��s�f��l�
B�O��`d��Pc7���,5�����s5���9���u"�k��C��.��Ww�ק�v��ė5n`�=���v�W�|�ͽ�Ý#b0���H�+��U@)bح�|�2hf&v����M%Oj�d6� ts9�a���b�Л_?T�]l*��� �dL��T%��	;���!��Qs�t�,v�]�ƢV�>�b���ǒI �7a��6��׮c��P���\���TQ �E$����;�d7hhn_yBXzr����p�-)�۝����aIN?/�"|B=W��[��hԉ.�!B/�*���� ��o�?W�����/�ONXg�`��\6�)�9R�������H��xi��&�M��$f�g�
�K~��������4\�#{}PlNq�ݪ���ⶶ�W	ċ���Ne���u�7�8J��5gAj}Y���i��`T@�h��E�K%*�B����IPy��RNP��1�g��?J>����徱�9�L�����W~j��}��ܯ��1�� <�	��Z�����*x ��rj�����v�Xt��e͉�n-��z&yl�B2��ۄ��k���#��x|��g95�h������^k��w�?X��7�j7�l?6�u�IPkdk��W�5E���^�H,xw�h#���G�?S7U��k"K{�Ή`~��~~6������*�n���>�YKp���X����`�ޖ�!����p1]j�-7( �X��;��qS��eA�[-Z��A�{-��6y<y�]�lu�H�7��U^u7@3�݉�	5����dp]e����!>�B��~$X*�Ui ��$$Tֵ�A4�:���xG��mn�'���0��X����;bYd�5��IZ��P���gB3�5j��9��}k�����Q"nJ�Y�ښ�}wd�Rgڞ�]�n����Ty<�z�B���gj�rS7
� �zq�%�3
Y$˵~�Fݧ�v���`�{͙�K��7��ޕ�E��	jI6&�`da��~,82z�d�J���e�ۊ���);&T-A1d->B�$P|"�?!{"q���&�Ѡ�5���`�$/�K����9��c 	6u������
��#���t�*1�n�Į0W��}|�iq Ul���[��C+d 3}VQ�=b	�oJ��p}�zu�ߍa�H6	�s��>�Z���D}�/f��g4��4��^����\Z�c8n�$J0.�>�����:�Ԇ�G&�p�f�t]��@2lZB�fy�����4߹j�=�rО�{k��;�o��
���F���=R��
�ĥ�%�=�Ώ��
�~���z�6��}�-�����4��Mx=��������)�ˉ���Q3y'"̦��j��ʐ�*�w�+�Ucf�34)���y���@5M�d�HԆ��Ax�dnŨ%�M��Z�����,��aB��T����9��0��[�lQjZ��.����(�g�O-�5 戾D�O%�S���T���,g,�.�m+�F=�Aj]�=LU��Q�A���ki8�w����-�H��|���[��]��5cI���]�?S���\��cȟg|Z:,@h�v�R�F����q�w������U�܌\&�E�Y*E�셪J$c�%�[H'9��1�X>+à�%�� ��-�-�(�ʠ� &�����}-Y� �V�m។ӗ�e#O���a2e9֪����SC)]�V�2}�����OūEsq�H8,��ڌ�<� �O�����D�[^�e {F��u�fVPL�D�y���>'�%~�ih�]��|�M�놠��L\3�8��! �>��;w��>�T�>���i�'th�J��RX����p�E�p x��'l�$3 ÑTқa�V�L�W7��\�_���m��d/�QsaF6��BS
q3�`6�e��Ю�_-6�e�r�v�G��^���M��lQI���l^)��m�{d�V�Z?�Y�F��W�ȷ�(ؘ����1��������T�D�P�2�Qo�<���a5�"��JYUԀ�%�q��n��3�>���_���JS��=I��uC�iR�x��~Ƭ���E?�,�~�n��N7GY]$c�*ؖأF�(?{��§���6 B��-���U�� �/do �q���e^jGM�o��%�>LD�J�g^`B�T4Nc�W�y���x%l�$�{��[���Oȴ����X�l�.�!�;��<6����W�-�[̾��a�f���6Y$�*ؖ��������n�:�,N|�th?�iLV�;��SQv���Ѻ
�D6�]�p4���4m�l�f�eLS���n��T�]�K��@�5��:���;�5�D��G�%�g{��:��|i��()��+�*(jɭ�(k=,F"2�YkI��b�}�_��E���1Z
��	�u�M�M��:y�e0�sr}+�:?{�u>k��J�w�TFؒ9u���K�����]�{�B�|]2��׶��8�
�+��H�m��7�o��gS\Ԓ� |�-�q2g?��ػ�c���v��@�G�WJ )Ě�V肞m����m�단i��J
�&7��1Lxz�2���co�x���ӓd_&����nX5�c�*��@)Q�K�����c���1����ds�����CSm��j}�K)�W��P�C6T� 뽼_��j�TӳT�|���B��5���Fg�39ծx�9s�(Ȱ����m��O�����6P����S�)�!F���q�����VxN��.Ը����*h3s,��T��2�����#%n%Ʌ��FA0�|�6b��0wV�<�9���Y76�~�>�l�pQ:�-O2s%��.���G
����C�&�׉m�O���>n�(M�Q�%�PO� �y��f�y$����m{7R�Ƙ���!���?����疛�w�t�y<}�FڏNg�7
�,]��-x� IGW���,Ʀ�ݷ�{%ihV���G�u�������w6x����+���/v��푉����YZ'����R�N�gYGB�����MC2��{��s�]m���.��K3�P��wQ��MM�P�3�Ǥj͉��=3'O1���f�{��4û�E1/+F%(>wz@PΧƦst���؝�VNZ��+�Vfͮ��0a�d���qc�ie��{9�~
\�
��{-E��V�{�A1�v�0>�H�1*ER�$�8�?\yφ?n�x)�ϰ�H2F����n�o�����߸����_|�&�K��I�=jcqW͇��&0*�`>@D��R�h�L�F�2gl�]��Q���� 䅠��� ������ɠ�y ���wGh8�
��C�O�Y8�"�Jxa}3~��Z�;�
q#(e`��1�E}6z�&( ����H��	�s���������q�lFTd	���7/����z���j�	!��نV�B@<|Y��.#���=J��Q|�����φ �r��l1g�~��g+� YR��!3K�+_H����-�6�e&W�����*\S�o��%.������M�;��q�C�]]�ǹ;�U�U��������/8`=����¨4[-)�8��Jc�� ]+T���0�,ܠc 7 Qt� �8�ĸ:7}X!zM�7d��PJ{�4�o�%sPPO����s���s�o�/�3���6aj���y��f�ޚ3ӡ�J7�Q����9��24A�6}��r3rCS4E�=��� �AaG�Á�}�  !F��t�*u�i��I�(�oj񸲚J�-�E�e�K�w�����R����f�|�G��j����@6;,��z�ص��)+��ڇAc�/*G�4��zz��U�|r{�p����W�5g��E�������π"�Ub�(���.3J3��N%~$����~��@�p�a?�9�� �� ��7Ӑ@6�"	��"s9s�����B?�+֒TB���O0����p>-������*�V��L4,�^�M�[s����A��ؠ`��s�X����T=o�y6/~�+F��s\QZ�1�c�ں?�5ҹ�S��l`��D��F�����H15�|d�*�a�+��$���rs��I��]�ð�w`z�<��x�$�l(�����\_�q�~\�� ��ޅ݅���1����ҁ��'Z�Y�]Ƅ<�'��1p��>�Ag��6ȱ�6tJ��0!�^��k�g����Wj*#��5�DQ?�75j?�җ�9hZ�7�* $��:̱`���'{#jZ�G3�|qq2��M�5��/���l�ϴu��P����x�-�t������F�)޽>�8�����J�a����p��[��vJ�Jd՗Ӓ%TiH˿����4��Qf