��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&��n?��1ů��> K�-� �&�T�Ek/ֆ�\�놭5�DꢘP���+L+X�4��J��#�0�8���������l��jT��+�(���������6�MC!D�;�m�퓊D@v_p��䙋ⲝ��C_�6�Ռ��#�� ���	RD�4D��畓7���vn�H���0���fX����4 �CS�C`{��;�L����li��� y+����FD�p"��]���y��R��K�({� .؜M�������	^5���ɋ��&���&�@*���
e�� �t+���
_6��O<��7f�M��u���m(MrN����z�jL���@T`��M3��c�uQ�Y���%�dD���,�~^���y@Ga��(����C����	��G�86�S$��ɳT�ز8���:r��/y�[ݦڍ#A�����i�&<nU��<[5)�Z�-Ĭv���0t���d���"_���:�'-��d��*��q����_d�y�N-��~";#��������Y��؆���	6ZJnԷW��έ$Y�K�?�4���L�w�Wmiɶ��Y�?jx#*�i���F�m�E����O6T>]i�_�9;�!(��kH7�OS��_��[-M�((��lO�s�$�g�x7`��ZV�E���F��,9�j	@���]}<�ahb5~ãdl&I^�	v����-�@�@���	��!��d��`j[Q��� r��;f�i�.�m+UH7��/OV��c��������l��i��M��*'��?���G� SK�M��H?�ç��q;��)��Rȩ�"@���r��Ml>8!�S��L��EgeH]�8��>]GR=&���C��i�Za�z�,�F��h�q��^���wT�a���%�9�n��?~SИſ~�mu�OlIv�4'sT���/a��^��9��*��G�Fh�DM�_��CN�<�_Pg��O5��}s�%��m�o߫R���X�Q?��dK�Z|:�=��yw9����i�������h]���M��\�mLu��t�@�nU�����R��^�:7�`��t���i�싛�>̳�.�7����
L�G��4�:�8ݾKcf����k5���:z�6����I%�[m����X��AT�Ϟ�̼���\�E�Bd���'�d^|Ō��Q0�������l�.0��L�j�7���vD�Fw=��u���R䑁zg2
��]m�c�	��u���Nfo�=��|p�z�bzĺ&Ǣ�z�A�+�Gof�N�4����;�ft�I����$���P��!�/]웷��|v|ZA`f��F( ̒�`�dMD����7��ݒ��%�(`�k͢#7{^Z��V�k�2�׳G~�B�.���x��!��5�%����#�8XU � RK+���nN�N/�ȝ�A����{��jӔ���l�3d������b���Š^�ն�|f��� �gQ��B�d�G���,�ܢ!�V��}[�R��F����������h�8e6=<�
CS�>gݡ�P1��,���kuW����A6��q>�me�.b��.����Zcv�6� 1�D��Í��o���D��WPG�v�=��n��&`�I~�,��Kk�-s!�D��F���#0��T�WG.�F�1�*�K<MI�IJ?��yL��]�?@�"k�H0�����-�^-Y�<��i8���/�X�[�l���:y �1/G�W����s>gH/����.'zXl�Εg�q���*�*�����ʊ�9��HF��YBg�0��g,5	�Z|X}	ۊ������}�.��C��gٸ4̺2�h��v$�$pn����65�OY�Ԑr�4��mH�Q�) �sMV�.�4�u;����/��`0����C�B���v�>�4��H�X�n��{�9𕏧�I@
�Q�zBv>ӕ��(�z�T��&�L��C��ڬ; O�!�Ă��"*�RUIB݆��4�i���a>�ط�ΦiO2��D-�/�&m�g�`B���G����(xWpA�`m ��4��%y*0�J�/K ����|��uWA�-�ß-tx���5���b��A�T(WO��4�B�mXTyߒ�*s_����j�N��'��)�а������^U�&s����$��͠����]4Y�	�4�̋���/�s=��K�_�Ű�TW�,~=�6���{P��Oj�Y�'�������'&$��Ed:
��S�ƴb�Ý��w�6oJW��pF�Y<`�� [Y�#uYgT��C/�L�:,���MU5�h#�>���w&����<
[�O
�a���ae�&�Ge���N��Ŷ5��x��U� ���C|j�N�luRH�F�0�K�$	h���"�Սg�8�DʤX%��g��$�\� ;=�}|�����X!���F�ٸ0-�����L�6�`�������P��V��k�� �5�.Q U�V�+�v�K8��T���~VvD�w��R���ގ��ɕ�|N�;�M�iMevt�@���L�� I��<�#�U�]�5M�	�K�V�K�O��F��e���0����A*��������s�1c�U������b����_F㭛����R?�� [�,��YA�sn+�}Ov�g��u�bw��k�MW�B�6����t�k*l�D�$ M[Z!x��P�!
��Vڈ������`�	:u�6���LId��p`�Z>�#т�j���j�3�}����:�� ��j¯����h�Ai׿���
�Q��^e:8�����l𒃧i0�a#��.u���jVyA��������'bEEӑqd�C��%D��n̚G�9�z�����O���5Y�͆萧�O�y����{���2QK�������F�6B|��Y8-/����m1�@
2��~�<��7V��<*V=�D�W�ƶYSO@xG$�����/�QQ���3)��^��X����k���j����}	9�ɩ�,� �u	�a��`r1b�uy��k����\}����"�c�"Nck^r]����j@[�����+�H\@u�J��-kv��
k�l����J��ɕ�����r9�@Ώh�m�'����&z��)$;isP�I��=�"��^S�ؑ��� 4�*j������hx�Vɲ~���<�$�|�����m��q����Ă�ȭftE	e���)6_9��W�Hu�Z[T�u��N�w��k�"{*���bZ#8��U��d�'�#9��2�MN�Ғ2>�;.�;�dC����/I���)Gc��v\��r�[�M���[�Q��,@N�7��|�@M� u_�[i�*���<��Rރ��.	�
ݺ+����uE��T{J��>=$�'2�\�&���H�>��Cr?������4/ӈl�6)� ������݊���]1�F�Jq���)�0���Н��Y\���%��m�?��rn��3v�����׻قz/T��}+t��V����.@A�\8��ep��M���^!X���8s�~,mg�������S���\�e��4 ��A�/o|�����/O�;�̊���Y��>����v��\e��fn�����s�l�Eʱ3{��d�gB���Y�����ȑ��xEK�Դ�CLB1��mS�gE�$��>f��HmɎJ�,A��g�}.0�;��(2+��i=����`Hg
����aw���ܫ��~��먑�q11 �E��a��F�"T������Q��Y9��$��	�0�{��k���Lo�?YK��t��sp٪7�%E�$��O��x�I��Vm������"ia�^����j߂lT�s�.�e�ZC��d�I��@Mo#�Ii΢��C�w�I�g[�X]n$5�.��P�N1���q����ɞ4mIK	���lu	X���z��F<��J�S�� څUrA�8��s'w�T���,b@b�ؒb0'`tY$���@�1��v�7+�Z"�ƛuNw~�*t�QUjk�A��Mm \���bͽ^���;ڸA�ٿ�Y����/�[���Ե��\��m��zZ�Ձ��17F�+���g7x��C�8ƣ�W����E*ǹo�������#����`'�:���<�l\��Ӹ�a1��)h�U��*S��oT@��m��K]�g�3���/�W��i���6rN0�>���|�}E�ϣ��9V�@�[��}��R/;�'O������?�&`�g���s�IO�oP�.�e�겸o�����[���W	�Q$k��-	xt#IQ}����>�� ��4��Q����&�Vl.��<oH��Q��<�i��)Ľ��?`��
9�mks���x}{�5��󟚛[��DE�:'�SE׆�;*��j�*�YR���=d�(� ��� V6e0w'<��2	�� �&d?��a�XA0S�z H�M=Y�De�&o �Z�n���<b�K�.�&�J�$}
Y=�<N��-�8�~y}�Ej`�4u��h���ם�,{,m=>�R
	�I�Ai3�b���pSWF�.�Z�f1�kA8��[�W�C�oSU��Ew�
4� �]5�*��qfV�]*�p��u�׮K���A�l���O�vz���܍��b9��5_�F��9�����R}�GS'��g��]nq��݋�#߀l�#�e�4�go�o���L(V�_j�M�-#Q����Ʒ�)��i�b������S�.�"�O�z��Δ;�{p������K�!�@hP`}ww��); G�[�\VJ�� J�a����@+G�cvoԤXgƽș�gwo��OAoW���X�A�QS�f�p��S�&j��	k���-����5!`�;��Kl�S��TL�D�3F<���J�3nrP|���;�*�U��l]�Y�@Q����Gϼز�M;Ȉ& q�5	ʴ�}`���u[o㯯l�i��ƨ����H�,����RX�C�:뛴��'h?����vl��߅�h�y�Y������Ԛ�3#����V��0�
)�Y�+������?�AF'�
�j��H4��*�ýV�}�Q|궢F��N��؉�.������,Nb�������Є�5)W���l��5�ӊ4���(c�kh�{�ZW}C�0{?�&���?G@���Ɛ+��VZv5�[�|BBf�B��~��V�W@�J�J:�/�R�� ��+��FP�g4���(�{���p��_�V�{���ѝ��UkՁ���降_��v�\S#Ms�-������n���YI���������&��0A���%�p�����]��%�=s�h��ޡpO�m-�kǖ�nJ��5�cዻOB����n�]Q�.�I����ܠ�l�f��I�ɘ��I��9����W0ݪg�<���2.�N��W�Pᑩ���N�\I��B�R�1�ڠ�_<��h� ��1�:a=;3�f����^f4ģ�Q�=��g%�'��`����W���E���$g�y��?���&ze��h�0Mo��w��2�YhZ+�29D\�����FdQ�y��ף��'>�\�DJ���"Co
�����@��B{��+�%�&�"�^_�����ɘ���n��q�Q��)�뤂���늢j�ʮ=����ۑm@���Oj{��	���x�IPi8x�EQ�;#�;�xN�Z',:�Aӵ�w��D���%v�_�"j)"���v���-�!�ʇ}�M9u~�x�Vަd8È��4��WѪZh�l�_�������T��WJ�Z�i�*�r�Zϧآ`��*<ww,��	�TוV��;I_��364f��1��M::�����>&�*@�c�H����GjG���G��s���נ�DB�%r�T����;����
�#�L�׆�p~T� b����)C��5�~If��
���r�
Y�6�=�:�zŊwϧ�+&�ۃ0�(� `����2�"}�e\���)���K��V1+ �Ǚ}g'��=��o�;�aD�L�� ���u���<��8�i$D�v�~{�I��� Ն�IQB��D�{e�R\����hz+!Dhj��	��b�	�̵[��E'��(�?�R_W��yjj7n|u��j+�
��Hz��7�W�)�"��ek�t$(���A�0�#M�G�z��-D&ԟp����"� *�~��?��T���O�n��/�\0������048�w~��v�3G��"2�1
�l2ȥ��`Nן��A����UEܔ�7�H��h[k6+��g�?<���2��C:w]��?�U>"��AX��t��^Fa�-� i