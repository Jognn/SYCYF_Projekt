��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&��n?��1ů��> K�-� �&�T�Ek/ֆ�\�놭5�DꢘP���+L+X�4��J��#�0�8���������l��jT��+�(���������6�MC!D�;�m�퓊D@v_p��䙋ⲝ��C_�6�Ռ��#�� ���	RD�4D��畓7���vn�H���0���fX����4 �CS�C`{��;�L����li��� y+����FD�p"��]���y��R��K�({� .؜M�������	^5���ɋ��&���&�@*���
e�� �t+���
_6��O<��7f�M��u���m(MrN����z�jL���@T`��M3��c�uQ�Y���%�dD���,�~^���y@Ga��(����C����	��G�86�S$��ɳT�ز8���:r��/y�[ݦڍ#A�����i�&<nU��<[5)�Z�-Ĭv���0t���d���"_���:�'-��d��*��q����_d�y�N-��~";#��������Y��؆���	6ZJnԷW��έ$Y�K�?�4���L�w�Wmiɶ��Y�?jx#*�i���F�m�E����O6T>]i�_�9;�!(��kH7�OS��_��[-M�((��lO�s�$�g�x7`��ZV�E���F��,9�j	@���]}<�ahb5~ãdl&I^�	v����-�@�@���	��!��d��`j[Q��� r��;f�i�.�m+UH7��/OV��c��������l��i��M��*'��?���G� SK���mkݛq�K� xwC�3���~���H��=�עR�>�קp�.f�Q�P�����=�26�|P]��i��Tsp�PY�2�����l�g}��:? ]�wr\ q9J���?�&j��D��:]�N�>eX}>u��n��s����⯀ۋWjݜ|�$��n�/�A���{p/D^��f�����w���6���6+	��f%>����%YE\�`X7���6�0�ߎ�}9)s�� [�ꒉ�Zi9�fV��B��࡚}r�&��5��~�����h����vX���S/�_���d/(ZZM�����H~ޯ�)��Ӵ|	������	P����� ��'�wa�)`Qϻ���U��\���>�W�+l *�M,
+���S�iŐM�{4���pq�=v�e������7�����Î,ߵ�(h`�pӦ*<l�^%;���T?�G��	�(���C:�K�Vo�d<9o��^ y�`֙����l7gAܧ���.楾߱4P�v�1A���w�D�~�z���d�iH�*��!u�4��t��C�e�D��d�P������6�,X��R�/���T����7t7_�f.�;@.r �$�eV&O�Q�������`���w��ww�M( �t���q��З@d��������m�tڂ{��,`���!��E䐞�u����#�Z�Q	�j��G�1p�)��
re,���'�	�	�5�ʄ��d\b!;��A�UdI���٥+��	)�t., oF�K����U޳7�*�����}"��ZW���N�{	6ֹM�PL�_e T+�XAs{��o���W"t��f[�������h �]۝��Z�/a]geQ�֎�ݰ���>-}�ӒV0L5ꐇ��?��P��4�ˤ���/���,�>_��+ȶ٤�|g�ЇF�w�G��$�u5��I7=�L�P��V%�J���Bf���v��U���%R�L�0Ѧ�x#�����y��;�}�dK��ނ���ڋ�P8'���c�ʺX���jе��5��E7����Z��9h~�U�*����+q�eI��z���<����$�u:8��%`l}-�NB()���(�J�_!��K��m/ 
+�.��w�喇�J@N���hb�h]뾔bQ�[���
o)����������Y<�d[A6�cI8�֎�D�\o��#�O+Jn�B,��@�\+��O�}� ��D��%| xہp9��j���8� �����濌gJ�G�%W�$�[��̺��y2�7hj1W�\���'�iR����)偫�O��e�I�E���Xe9�A�XV�c}�=�N�"^a�
������㽨�����:)��c!x��|��z@��6גs'��I7�q��u������P�[��0�G�P6�2��|�S���9E��h�:~[�,�s���~%��wf&�h>�5IL�p� �sd?�^��qm�-�vd~I��L���V݃�vT����A�g��h3<�Sl)��� �a���#GՑa4�u�l��ؘ�F� �$��p��mBY	���I�F4�o���zY��b�G�md�dhi*�Tԛ�.�<�� ]�n(kvP�$�*g]�/��s���ӱ�p��{�T,e	���^C7��,c�\!��(N�C�&��$���OVu�5�]�Eɱ���r�/����
��?��v�Z�c7B�W̏� j�-��w�m��wO2��꡼�E�V5������l���� M����[�^V޵-���k��\�HO��e���:<�)D�
��t��T���(J̃�gs#�ր�h[O��N8���C�_�6#xo��$]����U�QB,�-�EC:�`�3G�m�
f�:<�|2*�z)�"H�{�Ofua!�~T=r"9ڽ�;[7,=��T'��~eyWehH��^�ا�i3�)Hu�~���Ϯ!�q!l@��,;��i�\#��/:�O�J��̉,�2����	{�Q�L��-@9E��_&�e��l�,Ry����5�s��U}	=EM��:?�)�[�Xa�_r���9$����	Y�>i�?��f"�M��"@
I�A5)b�G�^���m��eT�2�H��ɓ����7��yN�����Xţ���e��Cr@�,���.݃I�� c9��p���x&4&�uGWc��%��zCY*��Z�X,]v�i싵�,�.��	�9�����-�@B]�xg�7��*�7=�i�I4ɭ٬���#���y��?l
�:?k��Pz��I��&vڌvW�zt{���!����;	� �����]ѳ� X����coq�������|Py���������|�-Ũ�<2�.��P(��#
:����e6�`��3#��r�_�=$IPt�j�ӵZ@�6Zv9�AFXO2_�,������4���)����ȍ"q�z�?`~yCM�8��ļ�q�����WBЏ��bׇB��c/ی��{�?�sJ�=�щ�T���0�E�#K����y��X�����1��Hr6E	W��¨�3߫���u,��Jz&���$���/W]DJ��N`Q0�U�~d��VЈN�"\ �O`e!�*�M���
���	l÷��" k��ft�Yw8 ���E
�����+��/�g��zD�bqu!��<l$E����R������3!�U��@�\1M��ҿ�q�No��<�?/�WqT���{T+/A�������r&9i�����X�Zk*;�mF?Y��m�(ă;��zdDQ�<^f�5���l�<�D��`;]!��	|)Cn �$��8m�g���Ȩ ��WtDW���x<�����D��@M��̎B<�x���MT����$yiu���Ҁ�SQ�� acB�g5fɣ��f�M���<�w �u n� ����Gx�C'����Fv�꓿=�o@R���Sʕ�P��(oC�f�q��r�98A�0х���3�M1�eW��y�'��VŨ݊1�Q���i���\�yJ=(%)7:���Q#ۥ��<g�m�� �+;t������+�s�,M�2P
!�n���#ܯ$����Z���S��j
IЮ"P-D�A�(0��i��oۿ���JC��7S �|9;k���9>D�䛬����S��/�h1ˮI�H*h�tаl������Q�N�8E�h�q؅XEF=�;^��.�;���q�~��$���=U�e]��N����s��V��ٵ��<����鄋�>m���\X�.�]�uy�U��Sy�4�Ʌ�h�I�W`�>7�B��}&�m6��i�8B�\{P����H��^�|���X,��'ˤ�_���nu��5i���C|�k3L��^?�#N*��8z�ۋ�:wQ�x�6(O��1��H�'�����a��0�qw��&M��؊�6����ð���$�哘!�̥:��cDfG���I	� %�f��������cU�qy�P����>}�nvhr���0P�U˰&�I�#�n�T���O�@����R�ʮ�U�Ղ��c֝��JB���z�4Q�m�&����&v9�םU�@�;��MA'7��-�h�kR0ln�Pd!Jm�/o :5㚭�c�<HT��wѮ7�%N��� ��\��I��G��+�T<��׶�]�@1�� v�?�j_- �4��L��+B�|�3���*��2���u�c���Xi�ZM��xuȐR4"6�9�P�tWtz�з�
W"�.)�-VH�h��Z9���q\?�����#%!���x��/�M���;�S%kT�q��!��|��|��A j��\
t�C>Bʋ�X��/�c��K��t��U�N{UK8����+ӜAr��'����^=�<	4B���$�Kr79q�5�����s{�=�9)t����3hfC��F�6�����}j��mR꟎='*�&;�ƪE����� �0�.�2�J��z�#*��S���9�»L�U��s/0�,��^;VJ5"��y}lV��_,����j�㪟 �ӯ��:�Q
"��zk	7߾�S�ޡ�z�۴*ܿ#�8�'�KN$�Ó��;�1�#jw��{���"O�3V�vGVܜ��9���HQ�T�&Մ+��_����'������C�ŝ�õ襔�h��^[��D�̠�K�#�Qg��ɸ��pAM�͹c���
I��"��+s?�y
���Uq��v/Ʌ�$g�1�*�[��I��LX�N�<}���K�,�Y>nU��0�9���F>0�M�Ç)��w�צ8)+V��$0+�3�T�(�[R��4���c����������B~��uۛ��f�E��/��,+W�vP4�6���-�$��C�ᰓ�_NX駽"s!i![��r�����3��;�h1	��\�4j��+L�ؼ/CI8�Om��uE��c���j���M%�UpZ}��߾pn[x�x����1�Y&H߶����Qk̫����̇�/yRPѐb�kHb��M��Ok��C��l8�4b�[���N�b�9TA��Ij�vfXe��6�Z�WD��q�C�(�!���ߛ���B�i�
��uR���&��n��ë��ïw��rړxj£�	x�ȉkMzsMс��k��~iW�������PN!U�jG���ɨ�"���9��P} \�E�2������FW��v����@7�Y�F�̸�3{n��_M%�up�$�3!��[�Jmد�9&��\|��ͦ���_�Y�6��q���ڔ�{�[��k�o�!і��+��A�ϐ��7mt.;��%/ڢ���[nhj��`s0�IAq6�D�Ʊ_\��'��Md_Y�=8G���a��]BB_�	�$�A�`�ٱ2����[T8���FZ3u1�H@a�aZV�͕
d7@\/e�vjȻ, Lw��w�����=;�U��8.E����^ӯ뾃�?CR�;�����,[5Y��M縆��p��J�*:sD���4|���dQ�NN~����{<aOqW�C� �D�`�N2�s��qDޠ�!u��S�2#1g<������6��6@��U���l���b�P�VC� P>��;G*�)�� k���-�
�ص�&��?��!����0Dp	itH��䭇�=�����ՓNEv��
S!�ԊVX��=}�L��o���ޒIꏍa�N�G-��X�\1=R
�/}��9B�È���|G���$̒\�8�UoiN�_F�|;���%|v݀�y��]�_N2$#z5!֚oTqi=+q~F��+�|VK��q�L�8k{� ���W����;ww��#�kX;����PjC�|�=Jbd�e�kx��W�Պ��Sf�,�ف��"r~>�& 8�����ѥ�������ħK��7��j9��0)^>E��8'y���I��2T��4!E��\�ɗ�R���=�LQD!�WV�0����gh5����p�[rA�`W�VK0Ӯ�gC��q��t�9�ȇ�̫�;\7/�F���l�rlHI\�D֗�5:�Q�6��dX�� 6z���Q�\�}�[���;_�`l�j��9C���k��]�V�!)�[�4A�<�K?�z�f9�O^��2�k�:۹]�F��7������3��,�vT�g���P��vo���y�.`bç�X'%�Π����w�g3�g�ۊ|'������5���x� ޞ�τnŲ�%���ݽ��-q9C�%��\Ĩ�vl\�Ays���#���=!� ��g�5q�l�-הЍ{;�FO��2�f|m�?=}k1�Sk^sl&�I�D<�
�=�����+�y/��t�Y�'��E�}�
�O��S���
*��)E4����d����6<�C/���hy���"���6���ӟ���E�7��M�s^6�i�9��;�؅��V�o�����E�U�����omu1fߑѷ�;e���ֺor,(�3�"�25G<�z��̖�7c�DQ�_��\����t�]u:��wot��U�u���0ӵ��*�������֢^�sV&0(׉��]���ܬ)ۙ�b`<�~��3F����K��:P�KN���a<m�{�_��=�=�'x�'��t�/��Z�����]��
��ia�S�hX�%�e��p;���C���H�H�$��5e|�?�v$*�s�XOX�w���������y�K�7��T}��Ss�g+>��G���oa�e"�fU���jf�����uJ>^8ް*.�{���:&x�u|'\S�1�8��V�;���֑�.ֵw�x��d�;7߹X�0g7��au}�ܼ���z����>h�7���b�|��^��̚S����Lֳ4�����l8���}�����8[а�*]!��������p}�V}A��į�����)<�����zA���t����]Zu"!��Z�ϐ/�G�:�R R�<���,��S�ȗ���Q{�^$*�V<��~G1o�����j�w������u�=���
͑���i�BU6_�%�-�#I�ǧ�����V~bL�m�ZJ�-��9/��h�EX?"(�h>훑?�,0e�N����r��^F)h�OٌA\f5�@M�� �p��-c٘��+:�yH��\�as���$g�r�K�b9��b~!*s�,_R�>�R]I�?"�#�����T>�~�=S[x�lL�z��Rs|�����O�L��)�_�rDݗv2�S�>�p-�9�����zf�DX�<2%pFՒ>�P��0g�)�I�;Kb��nP\)X =r�u\��#Ř+�5�v?�ɠ�j:(��.��L� q�P�)�B>y&,/PS��2��
�В��e#����j��u�N�������D�`To�����h�*�d������ހ/i����E[<�H�=Kg��ږ�Z �~��w�-��ɒI?�a���`��0ҒZ��M�A�T^�2�ڛ������m�ы0�i3�?� >�0�%���{HR����Z&�;ef��P+@ܶ h���ua5��%����d����:����t�w��~5]��t�T_�U]U=������.	�@���~�����?��8�/�~Ƽ2��G�@�`!+��Wk��r����bHn��-�~�+=1r1�<�tܺF���V_��
��F�{;�� �ږ����	��$�ٲ�e�8�M�	+,A^�.Fe��;��A��(3<���a��~3{d�U/�����v=�V#��6~��}ĸ�8k�v�+;�����U\sc����oBE#��֥���dI������p��w�ߵ<'H�(��A���=�T`�3���v�S��2�������Ep�?��ۖ�1�ƽt�9i���?E7l�HM.�C*:��n�5��C)�a����?���dY��=/�}^��W�J���9#vk�2'Ē�=��v�F���׎���d;�o��8�e�E?�}��q���Չ���-8�z�wM+Q�q[z;G�l^F��P�Z�{����笮N��!`���	��嬵���{[!����GV&�1hr)�0E)�����؁�{�/U7א��ǒ\Q.�w^��kV��[KA��KUJ3$��#������-P��W�wu��e~\Sʾ���!����c�K7�Z~�������Mz{�� l\�-ܸ����Z�OTFJ���2�J=��؍uQ;MXF��ն/p^���0u��3*��v�R�M�]* }�R&�DY��/L=��I��uJ.��):��Q`\��SD�pSd�0&��9�m�ĩ�G�œW�épx�!A�����#����u��@2k�}�6��S����$~�WW+)�+٤�S)�ܦ�p��%�yg�L�й��^�9���,>���׊���������f/*&A,X?Xζ�)��' �b����!
�~�Y�N�4�"�X�yB���ID�O���q���q�w��W��� u��&!F��9�&貊�����D�(w�����>�E��+�N݀L�pH	L+�+���H�x��Z�tqA�O!��#�vd�$�w��F��ux /��lҋ��v"YH��qĐ��yu���ҹf���Ϲ����=��	u"��$Ƈxp��&G"�Q%�#�C�$��y�t��`ؘ�/R��UwI�6�4b��ź��f��D�_�r�c2�a}��
 P�O#?�b��5�)�$b(�����/9��f� JH�Qhs��d����y��8 ��v�Kd�]�-�r6�Λᑌ��;�o"�8@<*�C��M�������E�I�^h�:YbǗ��G�O��/`�YF�]}�qj;V3��o:��JjK41�:����^h  �C�`�!�� co�v� �z�&��{������#����!̈���"�DX��Dt�n��s�P�lQz����0���c�w�=����� �-�r�(B)4�Nbww�Ǝ�����:BM��M������Q��L&l�쨸9� >پS�K嘸Dj����Y����mpZ�<�"в���L߱��'"��೭3�v���a>��(T*�1�{�~x��K�H���X���R��n��;��f�7qI���.���kyj��ݐS�?@�ɮ��<�� ��6#��J*��bKp?��Z�<�{х�3o\p �d�0:p��a�������Vg�|i M(rò��vWm(�4j42A�!R�C{��,����D�t�LDÄu��Q��Q�$�Y~7V�|�����$Gr.o_�]y���af���J�Qz��a�u�a��6���ap�P�୾���$�Y�5�h��\H���I��*�S¯�s|��#��|�����dzШ(�x���3�lF٩D3����f����ќt��&EDM�u;KA�R�@ �,;&H�z5�������f��!��%;��}��8����jb38���ʮM��"SĻ�9��#aq��A�B`�#`�rl����;���0�>���N�$p�ϡ��6�CJ�I�����'�cv��wH�kn��FQ#Յ��K���x��Aw�U���?8v}#��\ň�{����._O�vXm�f�w�q|�-�I����ٚ���]���S���5 v>��I�y$��~�?���N��7\b �c�v'�&ì�{�(,%�ZEژ�VYi�c���;�6G�[�Փ0�R�9zU���i7K�ԥ�kΗP�����V�Z#���I�oR=+��i��Dvh��Br�p&���v�D�ȅ�Q��j�-�gЇ��m_W���l��i4��[.!K,���<��b��GƤb֥4�L?	���;u^���Vs�7i��Y�$�Ha��+�(g��A�
'P__��j��f�҄pB�e���B�%m�Zlh_N�N�-yOK9aq�W&Dg_+��T:e.0o5��añPA�S�}����8n�z{���0`��>�^���>bm��J�1i�hۗ�b���n��]��l����d��"6�3L.�@�e�O;:��;"[[VR�(s��m�+�Ո�F�]%erޖ�S �f	�`�'��܀�oַb�GH�����aO��p03�/��]�`��4���m�)�9/�$ɍ2�ȚVn����=��~��x��߭��˩r��a	�����}y6l9�D�vbނ5��ХG���d�6T2��'�ӉpT��~�èu�@�.����t����P�;�@�l���~���Zn�Cf5�[ݾ������`�,X�#�8*�F��i?�R�I ��V������dI�&��uc�ܑL�u������!6�ڴ��cf.�>��0ø�n�s��D���8#7U$g,��g6�G�����U+��8���("`�W4F�Ҝ��f�C�+:�Y0����reC�P^��?bX!���۹�djωi���DSj�:�S��?�]O@(��3_��{)9�DvO��^�u�Ɇ�C
�Ѐ�=��5���+UBO�f*ȇ�M��z��r<�7��]�F?.&]?c`�(�hN��������Hk���l�A�ЏIZ%���UE)̡��(�7�I��f��� ��\�nǸ{������q����+�� ��S��������$�?�`�JF*l�_��~ o�[K�����P�	��UL_�۴�u�Hf����z�L\�S�٘-η��&O ��r��	��rGҞ�,��]�ɫq���U�k��h!l�s��|�0t��Utk�&��Pߕ�\)�[�g���<oY��ɇ��"\����@z�q2�0�l� ��^�C� V�=ר]����C�|�}�Y{C�	�����MM=��C����ͰA��T�~rи`�qU��G����-g!�%�*�@ؼv&�%�m�T@y������P�#��Yn ��=���ҴA�18Ym�jb�����>��g~4�)�b�U�����	�bN�;�n�L���x��6t�Aq�q�[�=����2�u���>UgV�R���40��} �����u���R��u�����F�%\��,p�l������9���MU<��ׂ�����L��k�pY���UDp�J���'*�gt61��u�;�B���Q�zScGY�9���n�%���Qr}��[�
����(8\��[��Ʃ���ٺ�IȬ�V�=��� ����D��@[%dk��/��ET�·P ����NP��՗��������f�3>��eS=0�K:�w��sv��*���>I��; �7{�j[aA/ug!3F���\��\��� ��g�!z9ՅL�O9@�ͧ�e������tD��w1��D �UR&)�gI"�&+:�`�Ms���=�-2��M�M�g��.���f=�ۺO9�C�E8��L�H�l��(y@�sk#hjG{Rf��D贅#ʘ��#`�v��I"��O���Ze��#x�v�^�n���iTgW�:�^��K�MK�-@���y�����U����3��G�9�(�|��2�#�������n�C��]%��1PĶ1c�#����YÁ�7��XB���+������rc�coW�W��u��,����<C`�*��/Tg3� �x���Њ�Q������Dj/��;�+�Ͽ����]I#�*�fv�F�D�!� 4Fy�*�y�~�_�ƪ�hˏ�2��eG<sUE��_zai��6�כ]��I��*6]��V�շ�}o�����5���hu�TL>�+���e�>�3��y��Zj�YR2�>�f!�񼏦���kPQ���v��G\�a������w�
e5���w�	S��;.��<�WF�#����1�}[t��1�F�J1��d9)�W���6HM��oɔ:�fS�0,,�G���s�<6�~q^��Hn��p� \^0?)��Q
��;�7��s��&�ǃ�mp�^!���FN�CE�z���}����>qU�1ǖ�9(�r��݁��9�E���O��O�6>Hm��b�Z���5D}g,��\�~����������]�ȷ�Þ���W"W�g;�g5����L? Ĥ�"����0~�|O�jw�7t˖Dbo�	�_n����_��
`r~��TJ�ro�id�>0,�}�-�Tt���������wL�����L.P�%u����4��mt��c�0���y���o�*��.\e`��9\б�8M?�\+�u����`�m	E �
<kbP����A]9���~?�)H����%s���_�u �ݙ�b�% WbȚs����ڜ|S�W�Ѱь�*z0��QTA��(m���.=�4�v~*k�ܰ��>�9�ˈa��H<�L�<��(>�x��B!ę�*�Mqܫ�x�a�]"���m���V�'Ȇ#\����kr��n�N�%�Rv�s��̡�e5Q�!l"JQ�"!�I��=�~��9�`����T��Ƃ	 ��M�s��?, �\�5����!il���:53H�~髮g&K����Q�W����bIp��u�[�I��R�~�4~�+�M[�h&�۸�k���$��~�!�w�+�6-D/z@E�	�S�}�hB��ǰx�Y_;��
��"�b
�Fv^�k�XoͶR���V�Ύ-��-�3��DC�RPW*!�՜	��o��X���y����O`����6�%�(���uz0�GU���K(>^NK��Q0�.������a:B�vM� ��;J�W�~�:�;n*K�Fg���+��#�H�-l����6�r��Z�-	�)����젻!�+^C�N��bgq��{ƿ����}�v������Me���C��.��iҌ!���� ��_��бf��- @k���5ND�ZLa̸�,�XвW�&�S<.�lŴHs�[1�ۙRG%5 z�����dP��,�~��)!/��aQ'[�����ɶ���T?��@k�/��q�<c	�X���82Y����xR_"e���m�W�|ޚa�I�lz�**I6���j�h���hq[U�)ޅ6������[�$!b���n�\���`��UF-�F�ɧ����*�Feih�m����ڍ�=B��n�*�ߚ=^Rg�S`��Q��7�t���}�$��l���(�b�U���
�;]b����ߒ���� �I��aT=l��2k8idz��a�	��EK8HޢJ�8y�I��b#8��~�N1����J�
������X�����:"ԑ��� eYgq�ms�8"�r��&�a��=*�F!D���i0�[�zB���.sv�x�2��x���_��̺�^>�4�������4b{	���Z��ģm���4AM�1�N��x�@�d�G{Gx�ѯ5��Y�8w�t[��@#�qT��!1��	¹���F#r.⅔�3��4��cQ}$ň��]KFY\>e�A���ײ0�!܁����琴7�k�Jd��jt@�2���Fg�[�P��bLn%���D]�|������_2x����O���}�K��t�$x�fdN�V���s�e$1������%Գ��1ܖ�hU3�Jg,@5n��-<��' �����ƀ�㢁�e���h*��j�!��9��Yэ¤��~TC�w0E�{��8v���D�(��g�H},�;����ؾ�^�9u>N�'J�ږ���v�~��;�c-YXP� �sߧ����h�}zA^ fR'� �ю�2LA�=���穨j�0���eb�CH�˞mH\b��Zt>�9[��	I�V�9�ꡞ�9������������KT���-gJ�@ɑ�ƽ������RG<:%�.؍�ߨ����I��B�>k����񲯾���΄K��銨�u�Xm�z��I~��&�b�Ij�{E��e�Nn+�D�Z#�Z��Њ�G�6~�[cl���s0�ðݜ���X��ηJp�[A󍢲�/���4N�oH��,���x q?�Xb��]#�S���½�8_�x���Ǖ�Ϸ�+����jp	D�v�*�_�n���}��Vtv�c6]^�A_+L�Y-CP+K��?ʾ�|����t"�#ˤz-�:ŵ���F7*���;�d#����ݤ���[t�f;�yE���E���62s�\z����$X�n*]u����.~#"�B�L�+��P�4)����5�<���H��V`����Y���9��(Y��KvG�W������Bd����|{�]�T*a�/�*%A�7���
�H�4�+3J`�Q����z�v������˟=�I}�b)�y@���9xL���]���F�'���O�f�:�y�gJG"���l�8�٧��E,�5(�m��&�Kc�߮T6�Ģr�p�^��l���t�P���
[4sb�����mA.-&۰t��1��������*U}��a�/�Tq�O�iB`� �r*$�A\�*[���0q����O%�Z�ԗ�M6v�W<x�0�y�M�3��ƚ�����x��70��u�1ep/�@�f8�(u�/
}J��֔b
͢L�;o����'�|�]%w�dE��:�91#Nw�	�h�ٚg���lb�%�9{@Ws��Z��P�b���� >�)I�ڏ��d������/��j�?	�}�1��6�����!WχQO�������d}�5���l�� �~�u�"}����H���$��f��~�70�������#�M=ԉ�����c1UN����Dg��OV�q�	݁ŞF��B�#n�5���;Һ>i
Y��a���M���꯻MĂ�Ek��H��Ԕ9H1
�\����<�a��X��C5�f���v�����$W��/t���ĠR������m�Z�����5̌;��9�����Z�����{Z#�8�t�J�X��Pg�»?QE}A�@%o�ψ�-Z�(�v��<��r��}}Ƹ���ZwC��uGmt=�bxm�(����{�J�r�ΑF�
�96Br��O�Ь�� �����=�����T����^:�):ye��}�P�Z�?'{*�U�?�b����͍s���z��i����0Y�&t��5��-}��~�{t	�l���8��H@�Rx���k#Fgu.�(Bj]�$���`<a���>m�o!�Z� #L춈�X�[�{:����ߍ���/���o^8��Ue�Q�ؠ5s��L?�����#�V_��k�ИC�?µ"�'>]s;�9����'CΩ�ϟt��3��|�\KG�|�R��1E�޲���ʱ��e1���b�f�v-�@LlT�V;���B{�7����x�X���
�;N��pW�걫��?����/Թ޼X� e�|�HDr���׍0�ؑ9�sg��S<�Di�lX0܌��$lcs,@���d��BGU�M��'nqLS`��8&�'cP	W0"���� ,���Ħ#4��<O��Y�5&�wʸ�.��W<u괚��Ī}XW	K����m�� �V�����.�E�UޟR�L0(3�P.�y�ιf��[g����t{�p ���~E�-c� �S����%��RQ.UcB���B$���j7�ѻ#��x�p�m.���əia���5��8��+
�������Y����������J���Ց7u������5���R�{jA�[T���˜`���=h�lۚ�b�UW�0����luT��%���}OAi�E��s�d�.�=�������a���V��*����y����5f�.٩��ʧ~���8���ob���+[��r�wvȾϰ�3'��8�ljvJ�@N�=�pV�����?�U�'G(�������ܵ����I����r
Sb������s��bA�/Ѭ�����[K���㇔M{����Q?�d�Tu"�ć�
�mS��2d
���������{��|�}`,*�iLZ�z{{�.�5�\����#���,IeB��ܜM�m
�1Wڱ�����A����=��K�L��Y'��G����9�u�K���P�8X�N�#h���?��u}�x!��Ay�S������u�bU7���m6�-�pM���wB^��s�\x��k
�]��q)7B��0Z� -��x<�:���"��&����Q+� 