��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&��n?��1ů��> K�-� �&�T�Ek/ֆ�\�놭5�DꢘP���+L+X�4��J��#�0�8���������l��jT��+�(���������6�MC!D�;�m�퓊D@v_p��䙋ⲝ��C_�6�Ռ��#�� ���	RD�4D��畓7���vn�H���0���fX����4 �CS�C`{��;�L����li��� y+����FD�p"��]���y��R��K�({� .؜M�������	^5���ɋ��&���&�@*���
e�� �t+���
_6��O<��7f�M��u���m(MrN����z�jL���@T`��M3��c�uQ�Y���%�dD���,�~^���y@Ga��(����C����	��G�86�S$��ɳT�ز8���:r��/y�[ݦڍ#A�����i�&<nU��<[5)�Z�-Ĭv���0t���d���"_���:�'-��d��*��q����_d�y�N-��~";#��������Y��؆���	6ZJnԷW��έ$Y�K�?�4���L�w�Wmiɶ��Y�?jx#*�i���F�m�E����O6T>]i�_�9;�!(��kH7�OS��_��[-M�((��lO�s�$�g�x7`��ZV�E���F��,9�j	@���]}<�ahb5~ãdl&I^�	v����-�@�@���	��!��d��`j[Q��� r��;f�i�.�m+UH7��/OV��c��������l��i��M��*'��?���G� SK�M��H?�מqT'J,@�����"��g��K�����%h�"7���ǵך��Q�W�n�!��A=�s�.�pq/��kt���q��x����}��3fP��1(cՂ�^��^QP��$3^ ���f&�x���IԸ�b7��$@�������}d��OcPR�|�g�&�?�����O�j�6K��K����]��x����Ñ�q�=΂�J��f�/Ar(+kd��s�~�S��ֳ������^�I�:�/\���;��)|I�'��?M��������3��+M�n\��lܫ'�������8���έ�[�q��Kg1���P��l�(�^��s9�*������*�,?t��o��
��m�fO���v�t..�1K�N�0&�!�ՓiJ��V��9X��/�:��)m����6�]2,,�b}�Z�X1�-K�$=�<�_[p��Q;=��g�hv�۫~pU�ߦ�j�ĝ�H��O��M�U�����N���!d�G��~�0�G���������jt���68bV*�˓�(�� w�_x4�p�_����È�L�^+������L�eP�Ԗ&���H�5Ŋ��1�{i��9�Fh����.2c�Ȝ��v`˂ꦞ!qw�4�SK�l�)��+f�I�Ӥ��i-��su�C~A���@��Q�p�����A�%��M.L	�M��#���8���l�sܖ^�J&������?Yp�I!��嫕5�ZcN$ir}���tX�6+���w{n�|3�`��� j�!h������"o�e����7Xu�m�/0��r�|��@�0�&�+hJ-�-1�QkC����5�I,���z������Or��#��g��K�O�V��"+��v1nO�=�a�����&5�
F/ɓ��yK����d���uxN�Si���%K�|����{��ar��y�W�K���6�1�7ɫR�����3(�sf�����,V�d��=/-�`,sd�_jqz�x�=��:.���^�I\S׹��gᖿ��F��&ֲJf�����xz���ң?Ôj��T���"��:B`��>dF_��LS*�L�_W���U���H�t^���`��v>r~����P��!�L��K���h;���k��$m��I
�t�E#�mx�$�A��ʌ�i��g�UK��A�,��	��Ө����)�)*�Ɣ��ۓ���W����	�i�ݘb��;���D�=�uA��^dߖ�L	��bu�6�`7�$*�E\}K�)VQ>�5]QP�����:O�z�ơƃv��{��/3��5�(
1�˝cd!����둿�6(�k����Q�"Bi\;S4_���&n\g�O?,��zF�oL�+1���-E�P;��OBL��``�M��T�t%�ԫc�R ��9�
)�.
���S���	^#���V�)4��1���z/�/I	�+����p���0!��(���:FIM��fx�a�R����1@��'�s�������~�5۠�eh���ӭ��)
u)��)KS�a4��������!�1�CXy�QM
tH��Y
4� �MwhU>J����^�o���{��y9���n2���L�z���j��,ܴZ��I�r.Ə9�{��1}��XS9����0�\\Վa�U���MҾ�A&}��L:.��������\5�l܈gp"�g�s!u ��	62��9YNa�N����z�;��Q�M��S�`��	y�ߏ�9��=T��x(#�;!UΝ�)P5	�8�,zі�����_��3�f��T��Q����
��[+��K�]�Zqb����5��w��7"���?]:�~��|���D���prs�Ֆ���V�3ϔT���w�;>(�-�ȷm�����6���VI����4��e+�ԇ _N0�5ޥ��aɮ����t�$ͦ�5�4RK�.�'�{Z����̤������)���qڈ��*^&|71�Lڐ�u=�����;�A�A�o�	�����S�a�%f���&1Ŧ�I������#\=���*(/���<�p�mΣ�\��w��1R&�_�;2�N\�M��8T���L� ����nt���p1�1��o�Y$��<6��*~x���=����ܻ��M���Nv!�vX��#�P��
��V �W�~C�KCK�j�Djt%&S�S�n1�S{"NV�s���&́M��x	�:抎e����q=y���p��d�cX��?S�lBB[n�]0�N��ʜJY/��XZ�iy�qm䚅�O���X��3��;�Y��.���@�������̞ǲNY��oh�?q �!A���l��$�ӽ�=fd�]�*?�G���gV�{uQ�F��x��Ok ��JT��,|�"G�NpM}P(A5������UmfR��宙��ȩ\fx;R+`�=�
��>f�@��\H|J��.Ć��Y&	�R�u�+�r��-�.��.lrU`���p��#�:���)���TY�i�����>ko�r�Ƿb�Z[���������0j�b�z��W���V����6n���вx�[����L�L���I���O�8����t�3K��C��d�:�x�H'�Qǔ^5����p�B���2$�h�S[0�!��7�f��7_�[�1�2�7�+�tkp�,��9&�Vq��k�F�\Wp�����Uؓ7+=$��ԅql�Ia�8ލϙ�ꣳ��\�p���͘��4b9S��F,��?,�����pn9�lJ�*go�Yx�×��QMU����&��wfH�%��S>3��`7��"��8������3k��U�>F��`��6����ì"��a)}PS;у�J*������$O�&8n�j�wA��\-��0�u��W>x��������*(Ewir��Ngj[5���fd��3g�z�#>y��a��1R=+������"��*����~.!���6��'�P��A��oƿڻYi�_5!������uYM�}�S:�����}�_<���J��3����=�=��Gx��2�D:�EW�g��x�M��}( n2�����dNg��<�r@Iz�յ2���_᥹�]��qUus��:P��.�\-�S�_��__?������_QMj��"����zq�Wk5g:宫�%�i��N��Й�שּׁ�!��s���v�����[��-��/�Q8h�sBk�OѶۜ�u����uQ�.������r����0��i���u�h��!o���s6�x�l!7yO�L�]��|��p��X�����d�}:�~������9f<����<�i�>���("1�U��ѵzm��CKq���d��r���D����SI	M,pPz�,�����_]���2�۷�|�&Ll�M~,ߛ0�*s���}��Тs�1��, �7_\
�; .��Ɂ!�<���ʪ� pS�3p�W�[��<*iHP�c4M���5�4���ݪ�x�+$#O�Y��XI�X�_;1����p��zB�	7Xm�z�IϺу�8>���3���6��m|�i�/
^;�Y`���>��#�(pz�	���X$.DM^���S5�2s��2��s�9���"b��� ڄx�
�_N�Cs׊�g?7�M.Ԇs��ܸ S�~���9VN4���R�솥���8��!�r���w�ߠ�6q1��Y0�u5���"���`+}�Lw�^"�d��EeQ�l�������M���m�_
m2��v Ǚ=��m,���6^' \Y�_��ƅ��cxZv���\����j��\�I�B�9���6���H���~�:��JF%�ZJu�����Q.�(i� ��0�]%�ض����-�������rs�G�)��:�"ѐj�Z ңH�d�V�h)0iw���r�"{��S�^tԾ��]���H�(�΅ncR֩�����{*QU�g�Y�ǁ�*]�Zdw��nU�)���/��e��'L-I���X��?H��_�up���	�i���v˓�P m��)�1�yC��Uz���Rʝy�A�W���쌫���z��O��Hb��{�]�֝O�Y�UM���w/(�[��[`����J���b@�xI|��(h"�^κB��ŝČZ9�u�?L��G��"^HX����I,w�5�qn£ўsz<�U|�$��b��V)�)�HB�]eH�U�ތh��<�P�3������I��1{悢&]$!S�j�����z�\�e�3�:�����)bQ��4`�bDp�i���"=��i���c/&�d����U<|���4���3�L�h���?�מ�Ɠy~��� 
�����~ ���qfP�ÍVX���"TN� ��:Cw;Z�ꨲ%�B&dG�����*�ݸD5A6�r��F��w	�{�N�r%X�Y֭����������t4���l|Qܗ�����^3�RhM��z���H�ޙ�@��DG߫|��T�"�Ũq�DZ�0�>Pɻ-x����Ŷ��M?��� r|�bZ��6�����C��!j�Z��F�1"	3Be�����@������Ս��pC��%zO�a=��Z+}PuD�BtM���_xc����1X��6�Í��'��+G�r%�������'+P�}"h29�~{�77讗�B��u�`��7ZQ Rr���J����,2���Ȣ>��	�~��rn��X`T�ԸC����Tw������evNo/4��R��d7�΃�;��:��G���v������p�ډi+ۣ�9�F��={~������p�d�������0lC�T�߸�������<8
#�mž��d�29���U�]v4��?1������k�qQcɓ��l�������ĎP��~�7�v���~��p�� D���E|���́rZ�J�?�'䖞�����z��גS�1�&D��������S��~�|��K�y��(;d>��/c�F���0������D�tJkXt/��ae6lo���!�g���vi���d���\�G[ț�0�����ܱ��sA��k�S���{g%NA DE[-�Cu^]� _>��J�;Jq԰�$7��j6��ٳQA2��*�gz,1�,�aN;1�V]���ʟD�Dl��
�
dy����kMG�0p~[ܢl��|}������d�{��vS��{X+�M}�n�@ �3�,��[(��[6 �$���H�M2�G;���E x�[��]Ћ��|g���f�o�,H�L���m�)oz��~r�E��Ñ�%L�dM����}?��S��V��4�{�QV|�����I��/8̳`��o<�3i���2k�Źɹg1����SJ�_<&,��u�r҂�VJ=��q��Y���뷨/�D���D�I;�p�����/�v��0R�1u/��m�ρ����z��l�K84/�R.����B�ݐ��\���"E��bF�UGE$�X�?��^7�O.���V�t�.�$���A\�0�o2��t�̲&D���!��� ��v��A±c��ꥃ��X|��)bM�p����SkIL��Em
9����N��^muW�t�/,��&M���>Ɍ�,a�K`a��F�"�bx�����S�ҕ'��mc$ޖ�P�D���,���8�Zf��z]�k,)�=D�[�|����oTdcY��T�Qb�AlƬP]���^JKjX�B�<�}
t��'9����E�?$IXs0�{�.�y]� ��dZâ>h��~h���~�0���O����Rlh{>�-):>	�a�^����_�0%���1؅l%K�Ò�S�t����W���L�gG)P'5Z�_m����r)шL�[6( �.�xwW��\T��^�� >��ުSOz�7�@��L�Vn���c��kGJN"�d��7�<)Nk�^C�i��>f�l����k_�sH!��9��bP�y�U������X�FEu�z
��CI�3-��)�8��H=����U(ئ�~;��0�����,�+�N'j�N�U���Z�r�,Ӡ-�b����m)a�T�h"J��r�l��k����Q���J���oy2O��U�t'�f�,O����D�xp���s4�t��I�0��ԛ3#���	ԆHg�O�
?[���R*j��E���#+�
R2�5�=��(�(^�W�5�{���WpD�$�Ч���ɣ@Οi���]5�l糷1J��ގ.����Er5��7�p�ђȎ�N�ֈO�)s�0�)Vbs�;���eaAp�~T/<�'��s�QX ���c!��0�FxˏI�%X�KT��/p�fLkTa����'��g��T�����$���(�,�"�g_ &��n��.� �WO�W��n����7w�6WF���FB{^\����qͩO�̎:k<t#h��fn\M[�C����R��	"�%�LVxZRtN���G���t��Ffsљ����
��g�2�i<{^44��J'��-ɪ�k���ޙ*��/4]�)�@�ov���2��%����yi�C�?=�>hr�c�h��0>t�c�Pn�5-�ÒF_j[�#>趝h@0�{��!p�еkj���2͚���+K�]���EQ7/��e
po���zhԪ:���z���j��X��rT���������)i�=�$v���5��=.��f�+���ib3���	���7p�7M7����gw����Ofo�j�%���`�	�S(��٭���PyhUs�[��#()P�VY
c���ޚډv⩱��ϩ�o���11�SF�W�X
���f�!�4�t�}�f��|�h�7�6 Y!p%s�g\��}g6�d��_�j`a%~ԙgA+�Oȟ}�'�1��:��S{�H��J��i�;��OˊqN����` �Xr0���'�"���] *����Y^m!󈰞`�8�!M�
������j̳;��?���f{�=$��#������ �WWx�?r�xz�pٔ��"s�镡�Îǐ���;va���
�?���G+ ��u��򚢶Hɩ>���ן����I��T��.�'��9�&먵L����s���y����ʋT/{��`�sAQ�]�� �+���)�pw^8�>���a�i��mV��tꅔ������j��~��:�t��<>#��D&