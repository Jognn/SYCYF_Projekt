��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&��n?��1ů��> K�-� �&�T�Ek/ֆ�\�놭5�DꢘP���+L+X�4��J��#�0�8���������l��jT��+�(���������6�MC!D�;�m�퓊D@v_p��䙋ⲝ��C_�6�Ռ��#�� ���	RD�4D��畓7���vn�H���0���fX����4 �CS�C`{��;�L����li��� y+����FD�p"��]���y��R��K�({� .؜M�������	^5���ɋ��&���&�@*���
e�� �t+���
_6��O<��7f�M��u���m(MrN����z�jL���@T`��M3��c�uQ�Y���%�dD���,�~^���y@Ga��(����C����	��G�86�S$��ɳT�ز8���:r��/y�[ݦڍ#A�����i�&<nU��<[5)�Z�-Ĭv���0t���d���"_���:�'-��d��*��q����_d�y�N-��~";#��������Y��؆���	6ZJnԷW��έ$Y�K�?�4���L�w�Wmiɶ��Y�?jx#*�i���F�m�E����O6T>]i�_�9;�!(��kH7�OS��_��[-M�((��lO�s�$�g�x7`��ZV�E���F��,9�j	@���]}<�ahb5~ãdl&I^�	v����-�@�@���	��!��d��`j[Q��� r��;f�i�.�m+UH7��/OV��c��������l��i��M��*'��?���G� SKٜ¬'�Wx�R�4{�ŲFRe����v2�	��t; i�k	�7
U�<���<�l�r�pV��$b����}/L��&�q��!�}��r�i�+׮+(s@�����K]>*D��E5�R�b�g�������y1��	ET��r'7�*��l<$�!�O��n���^��rnLzŉa�c9�=�m2�3�QG@/f�mwV�B�~��߽����_��of����S���#y~�B-k��JD�)���u�iKT!@��y�W:1�'���SZ�u=֣j�R��0{6�b�{���	��H� �(����{��ʶ��PL�`�X�
_�"ɁÊ��|Z�O�ܳ��U�iG�]f
������/�2��%C��
C���E��,C��0Y�U����P\���"��d�)�p߯zn�,�`}4r�7)�e$�&��ӄ�U�h�ZD\)5\}�N���3Zg�ִF���P�_�iK�:�3R�5�#bU%�fC�,�����>�X���@wI�U[��CQ2{/�*�����_g]��d��A]YX�L7�_2΂���uI�\'7-ڑ�#-G�mi���mR�xٱ�� f�A�%#�$�"�_ �Z�M���#t>&�ip1kc��������:_�~�?<M��a�a�e�KH>�����XKv���D�S�.��!��"���[_R$dI��1AGL��:�d�m�e�j�V(�1��r3�(C�V��N����Yk>!�kCZ���y=���չ�Ոꟻ���To$J��o	��JA ��C �#DX�صc:^�X�Eb?����J�R��n-�����&�7��R+�|��y1����h���Y����t]��b͜��o5��gE��3��o��l�{Ty���p��}l���L`m��T�c@FE4$1�����Cc-���:�S1p��V[L�L �19́gQ�͂/�<�Fj�ǜ�D��)rP%o*�l,O�d62}7U���dz��ع�h���z��y/���l�����8��9n�l@0���G����b�K�W��21*dg�q�c����@���j�#m�ŀۥ�O�P�:~�HȚuH ��c����
����:���Wd�C�Q:|�5�s�\P�ߔFiR��]n/��b��檗ۻ�|�,��
�wѻ<U,���+x�&Yݞ��]�5��WȺ�e�����X&�M�bo�f<�p�\�8,�k�}��]_�U�S6��I�Ba�(�bw�벑�M9��z��jV\iխ2zTD?��#ϖ��k�Iz�RQ�@t������u�?R�7X��,�=�Ĺh1�m�G.���d�H6>��������T����]z#S+�Е}ȒÀ��&��(|�����w�6�jV�*���4�|#���/㸓LZu�ZIW�s�G��
���)ow���t�[��Ì��^Qضh��+®`������n�U�I!���]��#�t����'�Z���+�2�(�js��)qȯ��K13@ػ�c(x�`|7��������K 죠�P�Hs�-?"?����{�������:���z�q#�u���W�;@8}�[kk'�&�[t��<my�_wK�YN%�����ﮕP/2D����-�5F��&+�����.��ߡ��͋YA��&�t1A��n8y����~���m�r��T5�W����#��Pr��i8�p[۶�ȱWv�v��s�2!��z
'��>�c�u�T��?�8?�<d���V|+�Z�9G�>�g)�u�k�O�������N|Hx�%��DZ4&t�����Lo��_�ѓ�*�����ឹzaи�D�H�D�y��D���7�C��ε��i�������s-䷧~��T��b$��V�  .��N�*܁]�'�IJЇ3��9�Ͱm�������5��w��BIl���O�$3�rxמ+V���T�|	���
+�`K���3K��Oׯ�_k�����^C<j��H��پ��䂈�'t�WO���<�vڱs�`�l%b6M����!Ȭ��w�MZ�����a �=WK��n����P����|]���̌��qu�>�Ԯs%k���g�0����)�w�Ŋп�-����)�����g�l�&�M���;垤�)5��{��S0-3tS�pB�8���`�_������O^Y�O|6S�G��)W@���s�i��������ܙ����!_�3����:����d5W�G�ж����Q��7�1B˰�#L"�%��1Z�Z���������Y@mC!�7�?+[�a��f�GQˀ�Mi�y�ig�GL�qEcI�(�u?��fCDe�S��0���Y����-���x��I/�u�cw���f�54Z�~����?��栨���n�M�%�Q8�E��5T����H�0�ow�\�@����cJ�f@"#2�bkߓ1!��4���T�C-j�MtpR�-媂5pguB�)�F���N#��iXw�U�HO���D�4)�I.v���=��z� ���� ���qL,�RAk�!����C]�'1����&�^쏺��:1��/gN��l�я�ܺ�-�K��7���1e��y(`�Lnt��u^�[���#�#�a߂J_�!ɍ�4`��P��e��_�J��b��;�9h�)�����
���� +���2>�E��6V_�إ��󘹻�"囥v��Խ�*��T�"��_>�@���������*�*�����mY3�y餕�I�S��wʩ�_D�uq{:����{�m����K�^����D�� �(�³S�q��Z���v��06l`j�M����!pӏ/r0��Έ��#*�_V�
E<m5����m�R�-2۷���!���_Xa�[���i�p �W	ۓP�V�ü�`��e�d��MZÉ�,��MA�L@�� �j���0 �%���v�����V�rS-��n{�S׾b�	3;'�e@v3sr�FQ���:N`�%Qj}?9xP�mx����RWr�ȃ0҅4���)�V�1�t�"T��6�&�ԕ�e1�(8o(h���öH��o�4ŝ�5.�d�ĭ��z
:���&7�j�X=�J+H3�m�0X��},_D��ܚ_����~�	�$e�w2u.�dz�{���ɪ�7�v|!��2�Ѵ��ߣ}$Ǚ���l��k.���s:�i��"\t�^b@��i'�A�0,XȒ���c;�Jf��|Z��π���[�v��Xk��d�L	��5)nfR�پK�0��~0q�r���M�E�f iO�d�;�p�A�R����[�c��~o��kO� _�|���8�!f�@�3KZ�е��&-�k����OL��ѹӚ������EN%��{e���FYF��M�